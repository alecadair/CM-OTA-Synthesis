MACRO NMOS_S_89651636_X2_Y9
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_89651636_X2_Y9 0 0 ;
  SIZE 3440 BY 54600 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 47620 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 4460 1860 51820 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 680 2290 53920 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 50905 ;
    LAYER M1 ;
      RECT 1165 51155 1415 52165 ;
    LAYER M1 ;
      RECT 1165 53255 1415 54265 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 735 47375 985 50905 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 1595 47375 1845 50905 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 50905 ;
    LAYER M1 ;
      RECT 2025 51155 2275 52165 ;
    LAYER M1 ;
      RECT 2025 53255 2275 54265 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2455 47375 2705 50905 ;
    LAYER M2 ;
      RECT 1120 280 2320 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 690 700 2750 980 ;
    LAYER M2 ;
      RECT 1120 6160 2320 6440 ;
    LAYER M2 ;
      RECT 1120 10360 2320 10640 ;
    LAYER M2 ;
      RECT 690 6580 2750 6860 ;
    LAYER M2 ;
      RECT 1120 12040 2320 12320 ;
    LAYER M2 ;
      RECT 1120 16240 2320 16520 ;
    LAYER M2 ;
      RECT 690 12460 2750 12740 ;
    LAYER M2 ;
      RECT 1120 17920 2320 18200 ;
    LAYER M2 ;
      RECT 1120 22120 2320 22400 ;
    LAYER M2 ;
      RECT 690 18340 2750 18620 ;
    LAYER M2 ;
      RECT 1120 23800 2320 24080 ;
    LAYER M2 ;
      RECT 1120 28000 2320 28280 ;
    LAYER M2 ;
      RECT 690 24220 2750 24500 ;
    LAYER M2 ;
      RECT 1120 29680 2320 29960 ;
    LAYER M2 ;
      RECT 1120 33880 2320 34160 ;
    LAYER M2 ;
      RECT 690 30100 2750 30380 ;
    LAYER M2 ;
      RECT 1120 35560 2320 35840 ;
    LAYER M2 ;
      RECT 1120 39760 2320 40040 ;
    LAYER M2 ;
      RECT 690 35980 2750 36260 ;
    LAYER M2 ;
      RECT 1120 41440 2320 41720 ;
    LAYER M2 ;
      RECT 1120 45640 2320 45920 ;
    LAYER M2 ;
      RECT 690 41860 2750 42140 ;
    LAYER M2 ;
      RECT 1120 47320 2320 47600 ;
    LAYER M2 ;
      RECT 1120 51520 2320 51800 ;
    LAYER M2 ;
      RECT 690 47740 2750 48020 ;
    LAYER M2 ;
      RECT 1120 53620 2320 53900 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47375 1375 47545 ;
    LAYER V1 ;
      RECT 1205 51575 1375 51745 ;
    LAYER V1 ;
      RECT 1205 53675 1375 53845 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47375 2235 47545 ;
    LAYER V1 ;
      RECT 2065 51575 2235 51745 ;
    LAYER V1 ;
      RECT 2065 53675 2235 53845 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 775 47795 945 47965 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 1635 47795 1805 47965 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 2495 47795 2665 47965 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 6225 1365 6375 ;
    LAYER V2 ;
      RECT 1215 12105 1365 12255 ;
    LAYER V2 ;
      RECT 1215 17985 1365 18135 ;
    LAYER V2 ;
      RECT 1215 23865 1365 24015 ;
    LAYER V2 ;
      RECT 1215 29745 1365 29895 ;
    LAYER V2 ;
      RECT 1215 35625 1365 35775 ;
    LAYER V2 ;
      RECT 1215 41505 1365 41655 ;
    LAYER V2 ;
      RECT 1215 47385 1365 47535 ;
    LAYER V2 ;
      RECT 1645 4545 1795 4695 ;
    LAYER V2 ;
      RECT 1645 10425 1795 10575 ;
    LAYER V2 ;
      RECT 1645 16305 1795 16455 ;
    LAYER V2 ;
      RECT 1645 22185 1795 22335 ;
    LAYER V2 ;
      RECT 1645 28065 1795 28215 ;
    LAYER V2 ;
      RECT 1645 33945 1795 34095 ;
    LAYER V2 ;
      RECT 1645 39825 1795 39975 ;
    LAYER V2 ;
      RECT 1645 45705 1795 45855 ;
    LAYER V2 ;
      RECT 1645 51585 1795 51735 ;
    LAYER V2 ;
      RECT 2075 765 2225 915 ;
    LAYER V2 ;
      RECT 2075 6645 2225 6795 ;
    LAYER V2 ;
      RECT 2075 12525 2225 12675 ;
    LAYER V2 ;
      RECT 2075 18405 2225 18555 ;
    LAYER V2 ;
      RECT 2075 24285 2225 24435 ;
    LAYER V2 ;
      RECT 2075 30165 2225 30315 ;
    LAYER V2 ;
      RECT 2075 36045 2225 36195 ;
    LAYER V2 ;
      RECT 2075 41925 2225 42075 ;
    LAYER V2 ;
      RECT 2075 47805 2225 47955 ;
    LAYER V2 ;
      RECT 2075 53685 2225 53835 ;
  END
END NMOS_S_89651636_X2_Y9
