MACRO NMOS_S_65192303_X12_Y8
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_65192303_X12_Y8 0 0 ;
  SIZE 12040 BY 48720 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5450 260 5730 41740 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5880 4460 6160 45940 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 6310 680 6590 48040 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 21505 ;
    LAYER M1 ;
      RECT 1165 21755 1415 22765 ;
    LAYER M1 ;
      RECT 1165 23855 1415 27385 ;
    LAYER M1 ;
      RECT 1165 27635 1415 28645 ;
    LAYER M1 ;
      RECT 1165 29735 1415 33265 ;
    LAYER M1 ;
      RECT 1165 33515 1415 34525 ;
    LAYER M1 ;
      RECT 1165 35615 1415 39145 ;
    LAYER M1 ;
      RECT 1165 39395 1415 40405 ;
    LAYER M1 ;
      RECT 1165 41495 1415 45025 ;
    LAYER M1 ;
      RECT 1165 45275 1415 46285 ;
    LAYER M1 ;
      RECT 1165 47375 1415 48385 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 735 17975 985 21505 ;
    LAYER M1 ;
      RECT 735 23855 985 27385 ;
    LAYER M1 ;
      RECT 735 29735 985 33265 ;
    LAYER M1 ;
      RECT 735 35615 985 39145 ;
    LAYER M1 ;
      RECT 735 41495 985 45025 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 1595 17975 1845 21505 ;
    LAYER M1 ;
      RECT 1595 23855 1845 27385 ;
    LAYER M1 ;
      RECT 1595 29735 1845 33265 ;
    LAYER M1 ;
      RECT 1595 35615 1845 39145 ;
    LAYER M1 ;
      RECT 1595 41495 1845 45025 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 21505 ;
    LAYER M1 ;
      RECT 2025 21755 2275 22765 ;
    LAYER M1 ;
      RECT 2025 23855 2275 27385 ;
    LAYER M1 ;
      RECT 2025 27635 2275 28645 ;
    LAYER M1 ;
      RECT 2025 29735 2275 33265 ;
    LAYER M1 ;
      RECT 2025 33515 2275 34525 ;
    LAYER M1 ;
      RECT 2025 35615 2275 39145 ;
    LAYER M1 ;
      RECT 2025 39395 2275 40405 ;
    LAYER M1 ;
      RECT 2025 41495 2275 45025 ;
    LAYER M1 ;
      RECT 2025 45275 2275 46285 ;
    LAYER M1 ;
      RECT 2025 47375 2275 48385 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2455 17975 2705 21505 ;
    LAYER M1 ;
      RECT 2455 23855 2705 27385 ;
    LAYER M1 ;
      RECT 2455 29735 2705 33265 ;
    LAYER M1 ;
      RECT 2455 35615 2705 39145 ;
    LAYER M1 ;
      RECT 2455 41495 2705 45025 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 21505 ;
    LAYER M1 ;
      RECT 2885 21755 3135 22765 ;
    LAYER M1 ;
      RECT 2885 23855 3135 27385 ;
    LAYER M1 ;
      RECT 2885 27635 3135 28645 ;
    LAYER M1 ;
      RECT 2885 29735 3135 33265 ;
    LAYER M1 ;
      RECT 2885 33515 3135 34525 ;
    LAYER M1 ;
      RECT 2885 35615 3135 39145 ;
    LAYER M1 ;
      RECT 2885 39395 3135 40405 ;
    LAYER M1 ;
      RECT 2885 41495 3135 45025 ;
    LAYER M1 ;
      RECT 2885 45275 3135 46285 ;
    LAYER M1 ;
      RECT 2885 47375 3135 48385 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3315 17975 3565 21505 ;
    LAYER M1 ;
      RECT 3315 23855 3565 27385 ;
    LAYER M1 ;
      RECT 3315 29735 3565 33265 ;
    LAYER M1 ;
      RECT 3315 35615 3565 39145 ;
    LAYER M1 ;
      RECT 3315 41495 3565 45025 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 21505 ;
    LAYER M1 ;
      RECT 3745 21755 3995 22765 ;
    LAYER M1 ;
      RECT 3745 23855 3995 27385 ;
    LAYER M1 ;
      RECT 3745 27635 3995 28645 ;
    LAYER M1 ;
      RECT 3745 29735 3995 33265 ;
    LAYER M1 ;
      RECT 3745 33515 3995 34525 ;
    LAYER M1 ;
      RECT 3745 35615 3995 39145 ;
    LAYER M1 ;
      RECT 3745 39395 3995 40405 ;
    LAYER M1 ;
      RECT 3745 41495 3995 45025 ;
    LAYER M1 ;
      RECT 3745 45275 3995 46285 ;
    LAYER M1 ;
      RECT 3745 47375 3995 48385 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4175 17975 4425 21505 ;
    LAYER M1 ;
      RECT 4175 23855 4425 27385 ;
    LAYER M1 ;
      RECT 4175 29735 4425 33265 ;
    LAYER M1 ;
      RECT 4175 35615 4425 39145 ;
    LAYER M1 ;
      RECT 4175 41495 4425 45025 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 21505 ;
    LAYER M1 ;
      RECT 4605 21755 4855 22765 ;
    LAYER M1 ;
      RECT 4605 23855 4855 27385 ;
    LAYER M1 ;
      RECT 4605 27635 4855 28645 ;
    LAYER M1 ;
      RECT 4605 29735 4855 33265 ;
    LAYER M1 ;
      RECT 4605 33515 4855 34525 ;
    LAYER M1 ;
      RECT 4605 35615 4855 39145 ;
    LAYER M1 ;
      RECT 4605 39395 4855 40405 ;
    LAYER M1 ;
      RECT 4605 41495 4855 45025 ;
    LAYER M1 ;
      RECT 4605 45275 4855 46285 ;
    LAYER M1 ;
      RECT 4605 47375 4855 48385 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5035 17975 5285 21505 ;
    LAYER M1 ;
      RECT 5035 23855 5285 27385 ;
    LAYER M1 ;
      RECT 5035 29735 5285 33265 ;
    LAYER M1 ;
      RECT 5035 35615 5285 39145 ;
    LAYER M1 ;
      RECT 5035 41495 5285 45025 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 21505 ;
    LAYER M1 ;
      RECT 5465 21755 5715 22765 ;
    LAYER M1 ;
      RECT 5465 23855 5715 27385 ;
    LAYER M1 ;
      RECT 5465 27635 5715 28645 ;
    LAYER M1 ;
      RECT 5465 29735 5715 33265 ;
    LAYER M1 ;
      RECT 5465 33515 5715 34525 ;
    LAYER M1 ;
      RECT 5465 35615 5715 39145 ;
    LAYER M1 ;
      RECT 5465 39395 5715 40405 ;
    LAYER M1 ;
      RECT 5465 41495 5715 45025 ;
    LAYER M1 ;
      RECT 5465 45275 5715 46285 ;
    LAYER M1 ;
      RECT 5465 47375 5715 48385 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 5895 17975 6145 21505 ;
    LAYER M1 ;
      RECT 5895 23855 6145 27385 ;
    LAYER M1 ;
      RECT 5895 29735 6145 33265 ;
    LAYER M1 ;
      RECT 5895 35615 6145 39145 ;
    LAYER M1 ;
      RECT 5895 41495 6145 45025 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 15625 ;
    LAYER M1 ;
      RECT 6325 15875 6575 16885 ;
    LAYER M1 ;
      RECT 6325 17975 6575 21505 ;
    LAYER M1 ;
      RECT 6325 21755 6575 22765 ;
    LAYER M1 ;
      RECT 6325 23855 6575 27385 ;
    LAYER M1 ;
      RECT 6325 27635 6575 28645 ;
    LAYER M1 ;
      RECT 6325 29735 6575 33265 ;
    LAYER M1 ;
      RECT 6325 33515 6575 34525 ;
    LAYER M1 ;
      RECT 6325 35615 6575 39145 ;
    LAYER M1 ;
      RECT 6325 39395 6575 40405 ;
    LAYER M1 ;
      RECT 6325 41495 6575 45025 ;
    LAYER M1 ;
      RECT 6325 45275 6575 46285 ;
    LAYER M1 ;
      RECT 6325 47375 6575 48385 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 6755 17975 7005 21505 ;
    LAYER M1 ;
      RECT 6755 23855 7005 27385 ;
    LAYER M1 ;
      RECT 6755 29735 7005 33265 ;
    LAYER M1 ;
      RECT 6755 35615 7005 39145 ;
    LAYER M1 ;
      RECT 6755 41495 7005 45025 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 15625 ;
    LAYER M1 ;
      RECT 7185 15875 7435 16885 ;
    LAYER M1 ;
      RECT 7185 17975 7435 21505 ;
    LAYER M1 ;
      RECT 7185 21755 7435 22765 ;
    LAYER M1 ;
      RECT 7185 23855 7435 27385 ;
    LAYER M1 ;
      RECT 7185 27635 7435 28645 ;
    LAYER M1 ;
      RECT 7185 29735 7435 33265 ;
    LAYER M1 ;
      RECT 7185 33515 7435 34525 ;
    LAYER M1 ;
      RECT 7185 35615 7435 39145 ;
    LAYER M1 ;
      RECT 7185 39395 7435 40405 ;
    LAYER M1 ;
      RECT 7185 41495 7435 45025 ;
    LAYER M1 ;
      RECT 7185 45275 7435 46285 ;
    LAYER M1 ;
      RECT 7185 47375 7435 48385 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M1 ;
      RECT 7615 17975 7865 21505 ;
    LAYER M1 ;
      RECT 7615 23855 7865 27385 ;
    LAYER M1 ;
      RECT 7615 29735 7865 33265 ;
    LAYER M1 ;
      RECT 7615 35615 7865 39145 ;
    LAYER M1 ;
      RECT 7615 41495 7865 45025 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 15625 ;
    LAYER M1 ;
      RECT 8045 15875 8295 16885 ;
    LAYER M1 ;
      RECT 8045 17975 8295 21505 ;
    LAYER M1 ;
      RECT 8045 21755 8295 22765 ;
    LAYER M1 ;
      RECT 8045 23855 8295 27385 ;
    LAYER M1 ;
      RECT 8045 27635 8295 28645 ;
    LAYER M1 ;
      RECT 8045 29735 8295 33265 ;
    LAYER M1 ;
      RECT 8045 33515 8295 34525 ;
    LAYER M1 ;
      RECT 8045 35615 8295 39145 ;
    LAYER M1 ;
      RECT 8045 39395 8295 40405 ;
    LAYER M1 ;
      RECT 8045 41495 8295 45025 ;
    LAYER M1 ;
      RECT 8045 45275 8295 46285 ;
    LAYER M1 ;
      RECT 8045 47375 8295 48385 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M1 ;
      RECT 8475 12095 8725 15625 ;
    LAYER M1 ;
      RECT 8475 17975 8725 21505 ;
    LAYER M1 ;
      RECT 8475 23855 8725 27385 ;
    LAYER M1 ;
      RECT 8475 29735 8725 33265 ;
    LAYER M1 ;
      RECT 8475 35615 8725 39145 ;
    LAYER M1 ;
      RECT 8475 41495 8725 45025 ;
    LAYER M1 ;
      RECT 8905 335 9155 3865 ;
    LAYER M1 ;
      RECT 8905 4115 9155 5125 ;
    LAYER M1 ;
      RECT 8905 6215 9155 9745 ;
    LAYER M1 ;
      RECT 8905 9995 9155 11005 ;
    LAYER M1 ;
      RECT 8905 12095 9155 15625 ;
    LAYER M1 ;
      RECT 8905 15875 9155 16885 ;
    LAYER M1 ;
      RECT 8905 17975 9155 21505 ;
    LAYER M1 ;
      RECT 8905 21755 9155 22765 ;
    LAYER M1 ;
      RECT 8905 23855 9155 27385 ;
    LAYER M1 ;
      RECT 8905 27635 9155 28645 ;
    LAYER M1 ;
      RECT 8905 29735 9155 33265 ;
    LAYER M1 ;
      RECT 8905 33515 9155 34525 ;
    LAYER M1 ;
      RECT 8905 35615 9155 39145 ;
    LAYER M1 ;
      RECT 8905 39395 9155 40405 ;
    LAYER M1 ;
      RECT 8905 41495 9155 45025 ;
    LAYER M1 ;
      RECT 8905 45275 9155 46285 ;
    LAYER M1 ;
      RECT 8905 47375 9155 48385 ;
    LAYER M1 ;
      RECT 9335 335 9585 3865 ;
    LAYER M1 ;
      RECT 9335 6215 9585 9745 ;
    LAYER M1 ;
      RECT 9335 12095 9585 15625 ;
    LAYER M1 ;
      RECT 9335 17975 9585 21505 ;
    LAYER M1 ;
      RECT 9335 23855 9585 27385 ;
    LAYER M1 ;
      RECT 9335 29735 9585 33265 ;
    LAYER M1 ;
      RECT 9335 35615 9585 39145 ;
    LAYER M1 ;
      RECT 9335 41495 9585 45025 ;
    LAYER M1 ;
      RECT 9765 335 10015 3865 ;
    LAYER M1 ;
      RECT 9765 4115 10015 5125 ;
    LAYER M1 ;
      RECT 9765 6215 10015 9745 ;
    LAYER M1 ;
      RECT 9765 9995 10015 11005 ;
    LAYER M1 ;
      RECT 9765 12095 10015 15625 ;
    LAYER M1 ;
      RECT 9765 15875 10015 16885 ;
    LAYER M1 ;
      RECT 9765 17975 10015 21505 ;
    LAYER M1 ;
      RECT 9765 21755 10015 22765 ;
    LAYER M1 ;
      RECT 9765 23855 10015 27385 ;
    LAYER M1 ;
      RECT 9765 27635 10015 28645 ;
    LAYER M1 ;
      RECT 9765 29735 10015 33265 ;
    LAYER M1 ;
      RECT 9765 33515 10015 34525 ;
    LAYER M1 ;
      RECT 9765 35615 10015 39145 ;
    LAYER M1 ;
      RECT 9765 39395 10015 40405 ;
    LAYER M1 ;
      RECT 9765 41495 10015 45025 ;
    LAYER M1 ;
      RECT 9765 45275 10015 46285 ;
    LAYER M1 ;
      RECT 9765 47375 10015 48385 ;
    LAYER M1 ;
      RECT 10195 335 10445 3865 ;
    LAYER M1 ;
      RECT 10195 6215 10445 9745 ;
    LAYER M1 ;
      RECT 10195 12095 10445 15625 ;
    LAYER M1 ;
      RECT 10195 17975 10445 21505 ;
    LAYER M1 ;
      RECT 10195 23855 10445 27385 ;
    LAYER M1 ;
      RECT 10195 29735 10445 33265 ;
    LAYER M1 ;
      RECT 10195 35615 10445 39145 ;
    LAYER M1 ;
      RECT 10195 41495 10445 45025 ;
    LAYER M1 ;
      RECT 10625 335 10875 3865 ;
    LAYER M1 ;
      RECT 10625 4115 10875 5125 ;
    LAYER M1 ;
      RECT 10625 6215 10875 9745 ;
    LAYER M1 ;
      RECT 10625 9995 10875 11005 ;
    LAYER M1 ;
      RECT 10625 12095 10875 15625 ;
    LAYER M1 ;
      RECT 10625 15875 10875 16885 ;
    LAYER M1 ;
      RECT 10625 17975 10875 21505 ;
    LAYER M1 ;
      RECT 10625 21755 10875 22765 ;
    LAYER M1 ;
      RECT 10625 23855 10875 27385 ;
    LAYER M1 ;
      RECT 10625 27635 10875 28645 ;
    LAYER M1 ;
      RECT 10625 29735 10875 33265 ;
    LAYER M1 ;
      RECT 10625 33515 10875 34525 ;
    LAYER M1 ;
      RECT 10625 35615 10875 39145 ;
    LAYER M1 ;
      RECT 10625 39395 10875 40405 ;
    LAYER M1 ;
      RECT 10625 41495 10875 45025 ;
    LAYER M1 ;
      RECT 10625 45275 10875 46285 ;
    LAYER M1 ;
      RECT 10625 47375 10875 48385 ;
    LAYER M1 ;
      RECT 11055 335 11305 3865 ;
    LAYER M1 ;
      RECT 11055 6215 11305 9745 ;
    LAYER M1 ;
      RECT 11055 12095 11305 15625 ;
    LAYER M1 ;
      RECT 11055 17975 11305 21505 ;
    LAYER M1 ;
      RECT 11055 23855 11305 27385 ;
    LAYER M1 ;
      RECT 11055 29735 11305 33265 ;
    LAYER M1 ;
      RECT 11055 35615 11305 39145 ;
    LAYER M1 ;
      RECT 11055 41495 11305 45025 ;
    LAYER M2 ;
      RECT 1120 280 10920 560 ;
    LAYER M2 ;
      RECT 1120 4480 10920 4760 ;
    LAYER M2 ;
      RECT 690 700 11350 980 ;
    LAYER M2 ;
      RECT 1120 6160 10920 6440 ;
    LAYER M2 ;
      RECT 1120 10360 10920 10640 ;
    LAYER M2 ;
      RECT 690 6580 11350 6860 ;
    LAYER M2 ;
      RECT 1120 12040 10920 12320 ;
    LAYER M2 ;
      RECT 1120 16240 10920 16520 ;
    LAYER M2 ;
      RECT 690 12460 11350 12740 ;
    LAYER M2 ;
      RECT 1120 17920 10920 18200 ;
    LAYER M2 ;
      RECT 1120 22120 10920 22400 ;
    LAYER M2 ;
      RECT 690 18340 11350 18620 ;
    LAYER M2 ;
      RECT 1120 23800 10920 24080 ;
    LAYER M2 ;
      RECT 1120 28000 10920 28280 ;
    LAYER M2 ;
      RECT 690 24220 11350 24500 ;
    LAYER M2 ;
      RECT 1120 29680 10920 29960 ;
    LAYER M2 ;
      RECT 1120 33880 10920 34160 ;
    LAYER M2 ;
      RECT 690 30100 11350 30380 ;
    LAYER M2 ;
      RECT 1120 35560 10920 35840 ;
    LAYER M2 ;
      RECT 1120 39760 10920 40040 ;
    LAYER M2 ;
      RECT 690 35980 11350 36260 ;
    LAYER M2 ;
      RECT 1120 41440 10920 41720 ;
    LAYER M2 ;
      RECT 1120 45640 10920 45920 ;
    LAYER M2 ;
      RECT 690 41860 11350 42140 ;
    LAYER M2 ;
      RECT 1120 47740 10920 48020 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 17975 1375 18145 ;
    LAYER V1 ;
      RECT 1205 22175 1375 22345 ;
    LAYER V1 ;
      RECT 1205 23855 1375 24025 ;
    LAYER V1 ;
      RECT 1205 28055 1375 28225 ;
    LAYER V1 ;
      RECT 1205 29735 1375 29905 ;
    LAYER V1 ;
      RECT 1205 33935 1375 34105 ;
    LAYER V1 ;
      RECT 1205 35615 1375 35785 ;
    LAYER V1 ;
      RECT 1205 39815 1375 39985 ;
    LAYER V1 ;
      RECT 1205 41495 1375 41665 ;
    LAYER V1 ;
      RECT 1205 45695 1375 45865 ;
    LAYER V1 ;
      RECT 1205 47795 1375 47965 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 17975 2235 18145 ;
    LAYER V1 ;
      RECT 2065 22175 2235 22345 ;
    LAYER V1 ;
      RECT 2065 23855 2235 24025 ;
    LAYER V1 ;
      RECT 2065 28055 2235 28225 ;
    LAYER V1 ;
      RECT 2065 29735 2235 29905 ;
    LAYER V1 ;
      RECT 2065 33935 2235 34105 ;
    LAYER V1 ;
      RECT 2065 35615 2235 35785 ;
    LAYER V1 ;
      RECT 2065 39815 2235 39985 ;
    LAYER V1 ;
      RECT 2065 41495 2235 41665 ;
    LAYER V1 ;
      RECT 2065 45695 2235 45865 ;
    LAYER V1 ;
      RECT 2065 47795 2235 47965 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 17975 3095 18145 ;
    LAYER V1 ;
      RECT 2925 22175 3095 22345 ;
    LAYER V1 ;
      RECT 2925 23855 3095 24025 ;
    LAYER V1 ;
      RECT 2925 28055 3095 28225 ;
    LAYER V1 ;
      RECT 2925 29735 3095 29905 ;
    LAYER V1 ;
      RECT 2925 33935 3095 34105 ;
    LAYER V1 ;
      RECT 2925 35615 3095 35785 ;
    LAYER V1 ;
      RECT 2925 39815 3095 39985 ;
    LAYER V1 ;
      RECT 2925 41495 3095 41665 ;
    LAYER V1 ;
      RECT 2925 45695 3095 45865 ;
    LAYER V1 ;
      RECT 2925 47795 3095 47965 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 17975 3955 18145 ;
    LAYER V1 ;
      RECT 3785 22175 3955 22345 ;
    LAYER V1 ;
      RECT 3785 23855 3955 24025 ;
    LAYER V1 ;
      RECT 3785 28055 3955 28225 ;
    LAYER V1 ;
      RECT 3785 29735 3955 29905 ;
    LAYER V1 ;
      RECT 3785 33935 3955 34105 ;
    LAYER V1 ;
      RECT 3785 35615 3955 35785 ;
    LAYER V1 ;
      RECT 3785 39815 3955 39985 ;
    LAYER V1 ;
      RECT 3785 41495 3955 41665 ;
    LAYER V1 ;
      RECT 3785 45695 3955 45865 ;
    LAYER V1 ;
      RECT 3785 47795 3955 47965 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 17975 4815 18145 ;
    LAYER V1 ;
      RECT 4645 22175 4815 22345 ;
    LAYER V1 ;
      RECT 4645 23855 4815 24025 ;
    LAYER V1 ;
      RECT 4645 28055 4815 28225 ;
    LAYER V1 ;
      RECT 4645 29735 4815 29905 ;
    LAYER V1 ;
      RECT 4645 33935 4815 34105 ;
    LAYER V1 ;
      RECT 4645 35615 4815 35785 ;
    LAYER V1 ;
      RECT 4645 39815 4815 39985 ;
    LAYER V1 ;
      RECT 4645 41495 4815 41665 ;
    LAYER V1 ;
      RECT 4645 45695 4815 45865 ;
    LAYER V1 ;
      RECT 4645 47795 4815 47965 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 17975 5675 18145 ;
    LAYER V1 ;
      RECT 5505 22175 5675 22345 ;
    LAYER V1 ;
      RECT 5505 23855 5675 24025 ;
    LAYER V1 ;
      RECT 5505 28055 5675 28225 ;
    LAYER V1 ;
      RECT 5505 29735 5675 29905 ;
    LAYER V1 ;
      RECT 5505 33935 5675 34105 ;
    LAYER V1 ;
      RECT 5505 35615 5675 35785 ;
    LAYER V1 ;
      RECT 5505 39815 5675 39985 ;
    LAYER V1 ;
      RECT 5505 41495 5675 41665 ;
    LAYER V1 ;
      RECT 5505 45695 5675 45865 ;
    LAYER V1 ;
      RECT 5505 47795 5675 47965 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12095 6535 12265 ;
    LAYER V1 ;
      RECT 6365 16295 6535 16465 ;
    LAYER V1 ;
      RECT 6365 17975 6535 18145 ;
    LAYER V1 ;
      RECT 6365 22175 6535 22345 ;
    LAYER V1 ;
      RECT 6365 23855 6535 24025 ;
    LAYER V1 ;
      RECT 6365 28055 6535 28225 ;
    LAYER V1 ;
      RECT 6365 29735 6535 29905 ;
    LAYER V1 ;
      RECT 6365 33935 6535 34105 ;
    LAYER V1 ;
      RECT 6365 35615 6535 35785 ;
    LAYER V1 ;
      RECT 6365 39815 6535 39985 ;
    LAYER V1 ;
      RECT 6365 41495 6535 41665 ;
    LAYER V1 ;
      RECT 6365 45695 6535 45865 ;
    LAYER V1 ;
      RECT 6365 47795 6535 47965 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12095 7395 12265 ;
    LAYER V1 ;
      RECT 7225 16295 7395 16465 ;
    LAYER V1 ;
      RECT 7225 17975 7395 18145 ;
    LAYER V1 ;
      RECT 7225 22175 7395 22345 ;
    LAYER V1 ;
      RECT 7225 23855 7395 24025 ;
    LAYER V1 ;
      RECT 7225 28055 7395 28225 ;
    LAYER V1 ;
      RECT 7225 29735 7395 29905 ;
    LAYER V1 ;
      RECT 7225 33935 7395 34105 ;
    LAYER V1 ;
      RECT 7225 35615 7395 35785 ;
    LAYER V1 ;
      RECT 7225 39815 7395 39985 ;
    LAYER V1 ;
      RECT 7225 41495 7395 41665 ;
    LAYER V1 ;
      RECT 7225 45695 7395 45865 ;
    LAYER V1 ;
      RECT 7225 47795 7395 47965 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6215 8255 6385 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12095 8255 12265 ;
    LAYER V1 ;
      RECT 8085 16295 8255 16465 ;
    LAYER V1 ;
      RECT 8085 17975 8255 18145 ;
    LAYER V1 ;
      RECT 8085 22175 8255 22345 ;
    LAYER V1 ;
      RECT 8085 23855 8255 24025 ;
    LAYER V1 ;
      RECT 8085 28055 8255 28225 ;
    LAYER V1 ;
      RECT 8085 29735 8255 29905 ;
    LAYER V1 ;
      RECT 8085 33935 8255 34105 ;
    LAYER V1 ;
      RECT 8085 35615 8255 35785 ;
    LAYER V1 ;
      RECT 8085 39815 8255 39985 ;
    LAYER V1 ;
      RECT 8085 41495 8255 41665 ;
    LAYER V1 ;
      RECT 8085 45695 8255 45865 ;
    LAYER V1 ;
      RECT 8085 47795 8255 47965 ;
    LAYER V1 ;
      RECT 8945 335 9115 505 ;
    LAYER V1 ;
      RECT 8945 4535 9115 4705 ;
    LAYER V1 ;
      RECT 8945 6215 9115 6385 ;
    LAYER V1 ;
      RECT 8945 10415 9115 10585 ;
    LAYER V1 ;
      RECT 8945 12095 9115 12265 ;
    LAYER V1 ;
      RECT 8945 16295 9115 16465 ;
    LAYER V1 ;
      RECT 8945 17975 9115 18145 ;
    LAYER V1 ;
      RECT 8945 22175 9115 22345 ;
    LAYER V1 ;
      RECT 8945 23855 9115 24025 ;
    LAYER V1 ;
      RECT 8945 28055 9115 28225 ;
    LAYER V1 ;
      RECT 8945 29735 9115 29905 ;
    LAYER V1 ;
      RECT 8945 33935 9115 34105 ;
    LAYER V1 ;
      RECT 8945 35615 9115 35785 ;
    LAYER V1 ;
      RECT 8945 39815 9115 39985 ;
    LAYER V1 ;
      RECT 8945 41495 9115 41665 ;
    LAYER V1 ;
      RECT 8945 45695 9115 45865 ;
    LAYER V1 ;
      RECT 8945 47795 9115 47965 ;
    LAYER V1 ;
      RECT 9805 335 9975 505 ;
    LAYER V1 ;
      RECT 9805 4535 9975 4705 ;
    LAYER V1 ;
      RECT 9805 6215 9975 6385 ;
    LAYER V1 ;
      RECT 9805 10415 9975 10585 ;
    LAYER V1 ;
      RECT 9805 12095 9975 12265 ;
    LAYER V1 ;
      RECT 9805 16295 9975 16465 ;
    LAYER V1 ;
      RECT 9805 17975 9975 18145 ;
    LAYER V1 ;
      RECT 9805 22175 9975 22345 ;
    LAYER V1 ;
      RECT 9805 23855 9975 24025 ;
    LAYER V1 ;
      RECT 9805 28055 9975 28225 ;
    LAYER V1 ;
      RECT 9805 29735 9975 29905 ;
    LAYER V1 ;
      RECT 9805 33935 9975 34105 ;
    LAYER V1 ;
      RECT 9805 35615 9975 35785 ;
    LAYER V1 ;
      RECT 9805 39815 9975 39985 ;
    LAYER V1 ;
      RECT 9805 41495 9975 41665 ;
    LAYER V1 ;
      RECT 9805 45695 9975 45865 ;
    LAYER V1 ;
      RECT 9805 47795 9975 47965 ;
    LAYER V1 ;
      RECT 10665 335 10835 505 ;
    LAYER V1 ;
      RECT 10665 4535 10835 4705 ;
    LAYER V1 ;
      RECT 10665 6215 10835 6385 ;
    LAYER V1 ;
      RECT 10665 10415 10835 10585 ;
    LAYER V1 ;
      RECT 10665 12095 10835 12265 ;
    LAYER V1 ;
      RECT 10665 16295 10835 16465 ;
    LAYER V1 ;
      RECT 10665 17975 10835 18145 ;
    LAYER V1 ;
      RECT 10665 22175 10835 22345 ;
    LAYER V1 ;
      RECT 10665 23855 10835 24025 ;
    LAYER V1 ;
      RECT 10665 28055 10835 28225 ;
    LAYER V1 ;
      RECT 10665 29735 10835 29905 ;
    LAYER V1 ;
      RECT 10665 33935 10835 34105 ;
    LAYER V1 ;
      RECT 10665 35615 10835 35785 ;
    LAYER V1 ;
      RECT 10665 39815 10835 39985 ;
    LAYER V1 ;
      RECT 10665 41495 10835 41665 ;
    LAYER V1 ;
      RECT 10665 45695 10835 45865 ;
    LAYER V1 ;
      RECT 10665 47795 10835 47965 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 775 18395 945 18565 ;
    LAYER V1 ;
      RECT 775 24275 945 24445 ;
    LAYER V1 ;
      RECT 775 30155 945 30325 ;
    LAYER V1 ;
      RECT 775 36035 945 36205 ;
    LAYER V1 ;
      RECT 775 41915 945 42085 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 1635 18395 1805 18565 ;
    LAYER V1 ;
      RECT 1635 24275 1805 24445 ;
    LAYER V1 ;
      RECT 1635 30155 1805 30325 ;
    LAYER V1 ;
      RECT 1635 36035 1805 36205 ;
    LAYER V1 ;
      RECT 1635 41915 1805 42085 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 2495 18395 2665 18565 ;
    LAYER V1 ;
      RECT 2495 24275 2665 24445 ;
    LAYER V1 ;
      RECT 2495 30155 2665 30325 ;
    LAYER V1 ;
      RECT 2495 36035 2665 36205 ;
    LAYER V1 ;
      RECT 2495 41915 2665 42085 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 3355 18395 3525 18565 ;
    LAYER V1 ;
      RECT 3355 24275 3525 24445 ;
    LAYER V1 ;
      RECT 3355 30155 3525 30325 ;
    LAYER V1 ;
      RECT 3355 36035 3525 36205 ;
    LAYER V1 ;
      RECT 3355 41915 3525 42085 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 4215 18395 4385 18565 ;
    LAYER V1 ;
      RECT 4215 24275 4385 24445 ;
    LAYER V1 ;
      RECT 4215 30155 4385 30325 ;
    LAYER V1 ;
      RECT 4215 36035 4385 36205 ;
    LAYER V1 ;
      RECT 4215 41915 4385 42085 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5075 18395 5245 18565 ;
    LAYER V1 ;
      RECT 5075 24275 5245 24445 ;
    LAYER V1 ;
      RECT 5075 30155 5245 30325 ;
    LAYER V1 ;
      RECT 5075 36035 5245 36205 ;
    LAYER V1 ;
      RECT 5075 41915 5245 42085 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 5935 18395 6105 18565 ;
    LAYER V1 ;
      RECT 5935 24275 6105 24445 ;
    LAYER V1 ;
      RECT 5935 30155 6105 30325 ;
    LAYER V1 ;
      RECT 5935 36035 6105 36205 ;
    LAYER V1 ;
      RECT 5935 41915 6105 42085 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 12515 6965 12685 ;
    LAYER V1 ;
      RECT 6795 18395 6965 18565 ;
    LAYER V1 ;
      RECT 6795 24275 6965 24445 ;
    LAYER V1 ;
      RECT 6795 30155 6965 30325 ;
    LAYER V1 ;
      RECT 6795 36035 6965 36205 ;
    LAYER V1 ;
      RECT 6795 41915 6965 42085 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 7655 12515 7825 12685 ;
    LAYER V1 ;
      RECT 7655 18395 7825 18565 ;
    LAYER V1 ;
      RECT 7655 24275 7825 24445 ;
    LAYER V1 ;
      RECT 7655 30155 7825 30325 ;
    LAYER V1 ;
      RECT 7655 36035 7825 36205 ;
    LAYER V1 ;
      RECT 7655 41915 7825 42085 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V1 ;
      RECT 8515 12515 8685 12685 ;
    LAYER V1 ;
      RECT 8515 18395 8685 18565 ;
    LAYER V1 ;
      RECT 8515 24275 8685 24445 ;
    LAYER V1 ;
      RECT 8515 30155 8685 30325 ;
    LAYER V1 ;
      RECT 8515 36035 8685 36205 ;
    LAYER V1 ;
      RECT 8515 41915 8685 42085 ;
    LAYER V1 ;
      RECT 9375 755 9545 925 ;
    LAYER V1 ;
      RECT 9375 6635 9545 6805 ;
    LAYER V1 ;
      RECT 9375 12515 9545 12685 ;
    LAYER V1 ;
      RECT 9375 18395 9545 18565 ;
    LAYER V1 ;
      RECT 9375 24275 9545 24445 ;
    LAYER V1 ;
      RECT 9375 30155 9545 30325 ;
    LAYER V1 ;
      RECT 9375 36035 9545 36205 ;
    LAYER V1 ;
      RECT 9375 41915 9545 42085 ;
    LAYER V1 ;
      RECT 10235 755 10405 925 ;
    LAYER V1 ;
      RECT 10235 6635 10405 6805 ;
    LAYER V1 ;
      RECT 10235 12515 10405 12685 ;
    LAYER V1 ;
      RECT 10235 18395 10405 18565 ;
    LAYER V1 ;
      RECT 10235 24275 10405 24445 ;
    LAYER V1 ;
      RECT 10235 30155 10405 30325 ;
    LAYER V1 ;
      RECT 10235 36035 10405 36205 ;
    LAYER V1 ;
      RECT 10235 41915 10405 42085 ;
    LAYER V1 ;
      RECT 11095 755 11265 925 ;
    LAYER V1 ;
      RECT 11095 6635 11265 6805 ;
    LAYER V1 ;
      RECT 11095 12515 11265 12685 ;
    LAYER V1 ;
      RECT 11095 18395 11265 18565 ;
    LAYER V1 ;
      RECT 11095 24275 11265 24445 ;
    LAYER V1 ;
      RECT 11095 30155 11265 30325 ;
    LAYER V1 ;
      RECT 11095 36035 11265 36205 ;
    LAYER V1 ;
      RECT 11095 41915 11265 42085 ;
    LAYER V2 ;
      RECT 5515 345 5665 495 ;
    LAYER V2 ;
      RECT 5515 6225 5665 6375 ;
    LAYER V2 ;
      RECT 5515 12105 5665 12255 ;
    LAYER V2 ;
      RECT 5515 17985 5665 18135 ;
    LAYER V2 ;
      RECT 5515 23865 5665 24015 ;
    LAYER V2 ;
      RECT 5515 29745 5665 29895 ;
    LAYER V2 ;
      RECT 5515 35625 5665 35775 ;
    LAYER V2 ;
      RECT 5515 41505 5665 41655 ;
    LAYER V2 ;
      RECT 5945 4545 6095 4695 ;
    LAYER V2 ;
      RECT 5945 10425 6095 10575 ;
    LAYER V2 ;
      RECT 5945 16305 6095 16455 ;
    LAYER V2 ;
      RECT 5945 22185 6095 22335 ;
    LAYER V2 ;
      RECT 5945 28065 6095 28215 ;
    LAYER V2 ;
      RECT 5945 33945 6095 34095 ;
    LAYER V2 ;
      RECT 5945 39825 6095 39975 ;
    LAYER V2 ;
      RECT 5945 45705 6095 45855 ;
    LAYER V2 ;
      RECT 6375 765 6525 915 ;
    LAYER V2 ;
      RECT 6375 6645 6525 6795 ;
    LAYER V2 ;
      RECT 6375 12525 6525 12675 ;
    LAYER V2 ;
      RECT 6375 18405 6525 18555 ;
    LAYER V2 ;
      RECT 6375 24285 6525 24435 ;
    LAYER V2 ;
      RECT 6375 30165 6525 30315 ;
    LAYER V2 ;
      RECT 6375 36045 6525 36195 ;
    LAYER V2 ;
      RECT 6375 41925 6525 42075 ;
    LAYER V2 ;
      RECT 6375 47805 6525 47955 ;
  END
END NMOS_S_65192303_X12_Y8
