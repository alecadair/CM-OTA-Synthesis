MACRO CURRENT_MIRROR_OTA
  ORIGIN 0 0 ;
  FOREIGN CURRENT_MIRROR_OTA 0 0 ;
  SIZE 13.02 BY 483.59 ;
  PIN ID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 2.87 2.78 3.15 32.5 ;
      LAYER M3 ;
        RECT 7.17 2.78 7.45 36.7 ;
      LAYER M3 ;
        RECT 2.87 18.715 3.15 19.085 ;
      LAYER M4 ;
        RECT 3.01 18.5 7.31 19.3 ;
      LAYER M3 ;
        RECT 7.17 18.715 7.45 19.085 ;
    END
  END ID
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 8.46 70.82 8.74 212.26 ;
      LAYER M3 ;
        RECT 6.74 64.1 7.02 476.02 ;
      LAYER M3 ;
        RECT 8.46 205.195 8.74 205.565 ;
      LAYER M4 ;
        RECT 6.88 204.98 8.6 205.78 ;
      LAYER M3 ;
        RECT 6.74 205.195 7.02 205.565 ;
    END
  END VOUT
  PIN VINN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 2.44 39.74 2.72 51.82 ;
    END
  END VINN
  PIN VINP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.6 39.74 7.88 51.82 ;
    END
  END VINP
  OBS 
  LAYER M3 ;
        RECT 1.58 70.82 1.86 212.26 ;
  LAYER M3 ;
        RECT 3.73 64.1 4.01 480.22 ;
  LAYER M3 ;
        RECT 6.31 68.3 6.59 480.22 ;
  LAYER M3 ;
        RECT 1.58 211.495 1.86 211.865 ;
  LAYER M4 ;
        RECT 1.72 211.28 3.87 212.08 ;
  LAYER M3 ;
        RECT 3.73 211.495 4.01 211.865 ;
  LAYER M4 ;
        RECT 3.87 211.28 6.45 212.08 ;
  LAYER M3 ;
        RECT 6.31 211.495 6.59 211.865 ;
  LAYER M3 ;
        RECT 1.58 211.495 1.86 211.865 ;
  LAYER M4 ;
        RECT 1.555 211.28 1.885 212.08 ;
  LAYER M3 ;
        RECT 3.73 211.495 4.01 211.865 ;
  LAYER M4 ;
        RECT 3.705 211.28 4.035 212.08 ;
  LAYER M3 ;
        RECT 1.58 211.495 1.86 211.865 ;
  LAYER M4 ;
        RECT 1.555 211.28 1.885 212.08 ;
  LAYER M3 ;
        RECT 3.73 211.495 4.01 211.865 ;
  LAYER M4 ;
        RECT 3.705 211.28 4.035 212.08 ;
  LAYER M3 ;
        RECT 1.58 211.495 1.86 211.865 ;
  LAYER M4 ;
        RECT 1.555 211.28 1.885 212.08 ;
  LAYER M3 ;
        RECT 3.73 211.495 4.01 211.865 ;
  LAYER M4 ;
        RECT 3.705 211.28 4.035 212.08 ;
  LAYER M3 ;
        RECT 6.31 211.495 6.59 211.865 ;
  LAYER M4 ;
        RECT 6.285 211.28 6.615 212.08 ;
  LAYER M3 ;
        RECT 1.58 211.495 1.86 211.865 ;
  LAYER M4 ;
        RECT 1.555 211.28 1.885 212.08 ;
  LAYER M3 ;
        RECT 3.73 211.495 4.01 211.865 ;
  LAYER M4 ;
        RECT 3.705 211.28 4.035 212.08 ;
  LAYER M3 ;
        RECT 6.31 211.495 6.59 211.865 ;
  LAYER M4 ;
        RECT 6.285 211.28 6.615 212.08 ;
  LAYER M3 ;
        RECT 2.01 43.94 2.29 56.02 ;
  LAYER M3 ;
        RECT 2.01 56.54 2.29 61.06 ;
  LAYER M3 ;
        RECT 1.15 66.62 1.43 208.06 ;
  LAYER M3 ;
        RECT 2.01 55.86 2.29 56.7 ;
  LAYER M3 ;
        RECT 2.01 60.9 2.29 66.78 ;
  LAYER M4 ;
        RECT 1.29 66.38 2.15 67.18 ;
  LAYER M3 ;
        RECT 1.15 66.595 1.43 66.965 ;
  LAYER M3 ;
        RECT 1.15 66.595 1.43 66.965 ;
  LAYER M4 ;
        RECT 1.125 66.38 1.455 67.18 ;
  LAYER M3 ;
        RECT 2.01 66.595 2.29 66.965 ;
  LAYER M4 ;
        RECT 1.985 66.38 2.315 67.18 ;
  LAYER M3 ;
        RECT 1.15 66.595 1.43 66.965 ;
  LAYER M4 ;
        RECT 1.125 66.38 1.455 67.18 ;
  LAYER M3 ;
        RECT 2.01 66.595 2.29 66.965 ;
  LAYER M4 ;
        RECT 1.985 66.38 2.315 67.18 ;
  LAYER M3 ;
        RECT 8.03 43.94 8.31 56.02 ;
  LAYER M3 ;
        RECT 8.03 56.54 8.31 61.06 ;
  LAYER M3 ;
        RECT 8.89 66.62 9.17 208.06 ;
  LAYER M3 ;
        RECT 8.03 55.86 8.31 56.7 ;
  LAYER M3 ;
        RECT 8.03 60.9 8.31 66.36 ;
  LAYER M2 ;
        RECT 8.17 66.22 9.03 66.5 ;
  LAYER M3 ;
        RECT 8.89 66.36 9.17 66.78 ;
  LAYER M2 ;
        RECT 8.01 66.22 8.33 66.5 ;
  LAYER M3 ;
        RECT 8.03 66.2 8.31 66.52 ;
  LAYER M2 ;
        RECT 8.87 66.22 9.19 66.5 ;
  LAYER M3 ;
        RECT 8.89 66.2 9.17 66.52 ;
  LAYER M2 ;
        RECT 8.01 66.22 8.33 66.5 ;
  LAYER M3 ;
        RECT 8.03 66.2 8.31 66.52 ;
  LAYER M2 ;
        RECT 8.87 66.22 9.19 66.5 ;
  LAYER M3 ;
        RECT 8.89 66.2 9.17 66.52 ;
  LAYER M3 ;
        RECT 3.3 6.98 3.58 36.7 ;
  LAYER M3 ;
        RECT 2.87 43.52 3.15 55.6 ;
  LAYER M3 ;
        RECT 7.17 43.52 7.45 55.6 ;
  LAYER M3 ;
        RECT 3.3 36.54 3.58 40.32 ;
  LAYER M2 ;
        RECT 3.01 40.18 3.44 40.46 ;
  LAYER M3 ;
        RECT 2.87 40.32 3.15 43.68 ;
  LAYER M3 ;
        RECT 2.87 43.915 3.15 44.285 ;
  LAYER M4 ;
        RECT 3.01 43.7 7.31 44.5 ;
  LAYER M3 ;
        RECT 7.17 43.915 7.45 44.285 ;
  LAYER M2 ;
        RECT 2.85 40.18 3.17 40.46 ;
  LAYER M3 ;
        RECT 2.87 40.16 3.15 40.48 ;
  LAYER M2 ;
        RECT 3.28 40.18 3.6 40.46 ;
  LAYER M3 ;
        RECT 3.3 40.16 3.58 40.48 ;
  LAYER M2 ;
        RECT 2.85 40.18 3.17 40.46 ;
  LAYER M3 ;
        RECT 2.87 40.16 3.15 40.48 ;
  LAYER M2 ;
        RECT 3.28 40.18 3.6 40.46 ;
  LAYER M3 ;
        RECT 3.3 40.16 3.58 40.48 ;
  LAYER M2 ;
        RECT 2.85 40.18 3.17 40.46 ;
  LAYER M3 ;
        RECT 2.87 40.16 3.15 40.48 ;
  LAYER M2 ;
        RECT 3.28 40.18 3.6 40.46 ;
  LAYER M3 ;
        RECT 3.3 40.16 3.58 40.48 ;
  LAYER M3 ;
        RECT 2.87 43.915 3.15 44.285 ;
  LAYER M4 ;
        RECT 2.845 43.7 3.175 44.5 ;
  LAYER M3 ;
        RECT 7.17 43.915 7.45 44.285 ;
  LAYER M4 ;
        RECT 7.145 43.7 7.475 44.5 ;
  LAYER M2 ;
        RECT 2.85 40.18 3.17 40.46 ;
  LAYER M3 ;
        RECT 2.87 40.16 3.15 40.48 ;
  LAYER M2 ;
        RECT 3.28 40.18 3.6 40.46 ;
  LAYER M3 ;
        RECT 3.3 40.16 3.58 40.48 ;
  LAYER M3 ;
        RECT 2.87 43.915 3.15 44.285 ;
  LAYER M4 ;
        RECT 2.845 43.7 3.175 44.5 ;
  LAYER M3 ;
        RECT 7.17 43.915 7.45 44.285 ;
  LAYER M4 ;
        RECT 7.145 43.7 7.475 44.5 ;
  LAYER M1 ;
        RECT 6.325 33.095 6.575 36.625 ;
  LAYER M1 ;
        RECT 6.325 31.835 6.575 32.845 ;
  LAYER M1 ;
        RECT 6.325 27.215 6.575 30.745 ;
  LAYER M1 ;
        RECT 6.325 25.955 6.575 26.965 ;
  LAYER M1 ;
        RECT 6.325 21.335 6.575 24.865 ;
  LAYER M1 ;
        RECT 6.325 20.075 6.575 21.085 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 18.985 ;
  LAYER M1 ;
        RECT 6.325 14.195 6.575 15.205 ;
  LAYER M1 ;
        RECT 6.325 9.575 6.575 13.105 ;
  LAYER M1 ;
        RECT 6.325 8.315 6.575 9.325 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 33.095 6.145 36.625 ;
  LAYER M1 ;
        RECT 5.895 27.215 6.145 30.745 ;
  LAYER M1 ;
        RECT 5.895 21.335 6.145 24.865 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 18.985 ;
  LAYER M1 ;
        RECT 5.895 9.575 6.145 13.105 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 33.095 7.005 36.625 ;
  LAYER M1 ;
        RECT 6.755 27.215 7.005 30.745 ;
  LAYER M1 ;
        RECT 6.755 21.335 7.005 24.865 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M1 ;
        RECT 6.755 9.575 7.005 13.105 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 33.095 7.435 36.625 ;
  LAYER M1 ;
        RECT 7.185 31.835 7.435 32.845 ;
  LAYER M1 ;
        RECT 7.185 27.215 7.435 30.745 ;
  LAYER M1 ;
        RECT 7.185 25.955 7.435 26.965 ;
  LAYER M1 ;
        RECT 7.185 21.335 7.435 24.865 ;
  LAYER M1 ;
        RECT 7.185 20.075 7.435 21.085 ;
  LAYER M1 ;
        RECT 7.185 15.455 7.435 18.985 ;
  LAYER M1 ;
        RECT 7.185 14.195 7.435 15.205 ;
  LAYER M1 ;
        RECT 7.185 9.575 7.435 13.105 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 9.325 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 33.095 7.865 36.625 ;
  LAYER M1 ;
        RECT 7.615 27.215 7.865 30.745 ;
  LAYER M1 ;
        RECT 7.615 21.335 7.865 24.865 ;
  LAYER M1 ;
        RECT 7.615 15.455 7.865 18.985 ;
  LAYER M1 ;
        RECT 7.615 9.575 7.865 13.105 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 33.095 8.295 36.625 ;
  LAYER M1 ;
        RECT 8.045 31.835 8.295 32.845 ;
  LAYER M1 ;
        RECT 8.045 27.215 8.295 30.745 ;
  LAYER M1 ;
        RECT 8.045 25.955 8.295 26.965 ;
  LAYER M1 ;
        RECT 8.045 21.335 8.295 24.865 ;
  LAYER M1 ;
        RECT 8.045 20.075 8.295 21.085 ;
  LAYER M1 ;
        RECT 8.045 15.455 8.295 18.985 ;
  LAYER M1 ;
        RECT 8.045 14.195 8.295 15.205 ;
  LAYER M1 ;
        RECT 8.045 9.575 8.295 13.105 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 9.325 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 33.095 8.725 36.625 ;
  LAYER M1 ;
        RECT 8.475 27.215 8.725 30.745 ;
  LAYER M1 ;
        RECT 8.475 21.335 8.725 24.865 ;
  LAYER M1 ;
        RECT 8.475 15.455 8.725 18.985 ;
  LAYER M1 ;
        RECT 8.475 9.575 8.725 13.105 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M2 ;
        RECT 6.28 36.4 8.34 36.68 ;
  LAYER M2 ;
        RECT 6.28 32.2 8.34 32.48 ;
  LAYER M2 ;
        RECT 5.85 35.98 8.77 36.26 ;
  LAYER M2 ;
        RECT 6.28 30.52 8.34 30.8 ;
  LAYER M2 ;
        RECT 6.28 26.32 8.34 26.6 ;
  LAYER M2 ;
        RECT 5.85 30.1 8.77 30.38 ;
  LAYER M2 ;
        RECT 6.28 24.64 8.34 24.92 ;
  LAYER M2 ;
        RECT 6.28 20.44 8.34 20.72 ;
  LAYER M2 ;
        RECT 5.85 24.22 8.77 24.5 ;
  LAYER M2 ;
        RECT 6.28 18.76 8.34 19.04 ;
  LAYER M2 ;
        RECT 6.28 14.56 8.34 14.84 ;
  LAYER M2 ;
        RECT 5.85 18.34 8.77 18.62 ;
  LAYER M2 ;
        RECT 6.28 12.88 8.34 13.16 ;
  LAYER M2 ;
        RECT 6.28 8.68 8.34 8.96 ;
  LAYER M2 ;
        RECT 5.85 12.46 8.77 12.74 ;
  LAYER M2 ;
        RECT 6.28 7 8.34 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 8.34 3.08 ;
  LAYER M2 ;
        RECT 5.85 6.58 8.77 6.86 ;
  LAYER M2 ;
        RECT 6.28 0.7 8.34 0.98 ;
  LAYER M3 ;
        RECT 7.17 2.78 7.45 36.7 ;
  LAYER M3 ;
        RECT 7.6 0.68 7.88 36.28 ;
  LAYER M1 ;
        RECT 3.745 64.175 3.995 67.705 ;
  LAYER M1 ;
        RECT 3.745 67.955 3.995 68.965 ;
  LAYER M1 ;
        RECT 3.745 70.055 3.995 73.585 ;
  LAYER M1 ;
        RECT 3.745 73.835 3.995 74.845 ;
  LAYER M1 ;
        RECT 3.745 75.935 3.995 79.465 ;
  LAYER M1 ;
        RECT 3.745 79.715 3.995 80.725 ;
  LAYER M1 ;
        RECT 3.745 81.815 3.995 85.345 ;
  LAYER M1 ;
        RECT 3.745 85.595 3.995 86.605 ;
  LAYER M1 ;
        RECT 3.745 87.695 3.995 91.225 ;
  LAYER M1 ;
        RECT 3.745 91.475 3.995 92.485 ;
  LAYER M1 ;
        RECT 3.745 93.575 3.995 97.105 ;
  LAYER M1 ;
        RECT 3.745 97.355 3.995 98.365 ;
  LAYER M1 ;
        RECT 3.745 99.455 3.995 102.985 ;
  LAYER M1 ;
        RECT 3.745 103.235 3.995 104.245 ;
  LAYER M1 ;
        RECT 3.745 105.335 3.995 108.865 ;
  LAYER M1 ;
        RECT 3.745 109.115 3.995 110.125 ;
  LAYER M1 ;
        RECT 3.745 111.215 3.995 114.745 ;
  LAYER M1 ;
        RECT 3.745 114.995 3.995 116.005 ;
  LAYER M1 ;
        RECT 3.745 117.095 3.995 120.625 ;
  LAYER M1 ;
        RECT 3.745 120.875 3.995 121.885 ;
  LAYER M1 ;
        RECT 3.745 122.975 3.995 126.505 ;
  LAYER M1 ;
        RECT 3.745 126.755 3.995 127.765 ;
  LAYER M1 ;
        RECT 3.745 128.855 3.995 132.385 ;
  LAYER M1 ;
        RECT 3.745 132.635 3.995 133.645 ;
  LAYER M1 ;
        RECT 3.745 134.735 3.995 138.265 ;
  LAYER M1 ;
        RECT 3.745 138.515 3.995 139.525 ;
  LAYER M1 ;
        RECT 3.745 140.615 3.995 144.145 ;
  LAYER M1 ;
        RECT 3.745 144.395 3.995 145.405 ;
  LAYER M1 ;
        RECT 3.745 146.495 3.995 150.025 ;
  LAYER M1 ;
        RECT 3.745 150.275 3.995 151.285 ;
  LAYER M1 ;
        RECT 3.745 152.375 3.995 155.905 ;
  LAYER M1 ;
        RECT 3.745 156.155 3.995 157.165 ;
  LAYER M1 ;
        RECT 3.745 158.255 3.995 161.785 ;
  LAYER M1 ;
        RECT 3.745 162.035 3.995 163.045 ;
  LAYER M1 ;
        RECT 3.745 164.135 3.995 167.665 ;
  LAYER M1 ;
        RECT 3.745 167.915 3.995 168.925 ;
  LAYER M1 ;
        RECT 3.745 170.015 3.995 173.545 ;
  LAYER M1 ;
        RECT 3.745 173.795 3.995 174.805 ;
  LAYER M1 ;
        RECT 3.745 175.895 3.995 179.425 ;
  LAYER M1 ;
        RECT 3.745 179.675 3.995 180.685 ;
  LAYER M1 ;
        RECT 3.745 181.775 3.995 185.305 ;
  LAYER M1 ;
        RECT 3.745 185.555 3.995 186.565 ;
  LAYER M1 ;
        RECT 3.745 187.655 3.995 191.185 ;
  LAYER M1 ;
        RECT 3.745 191.435 3.995 192.445 ;
  LAYER M1 ;
        RECT 3.745 193.535 3.995 197.065 ;
  LAYER M1 ;
        RECT 3.745 197.315 3.995 198.325 ;
  LAYER M1 ;
        RECT 3.745 199.415 3.995 202.945 ;
  LAYER M1 ;
        RECT 3.745 203.195 3.995 204.205 ;
  LAYER M1 ;
        RECT 3.745 205.295 3.995 208.825 ;
  LAYER M1 ;
        RECT 3.745 209.075 3.995 210.085 ;
  LAYER M1 ;
        RECT 3.745 211.175 3.995 214.705 ;
  LAYER M1 ;
        RECT 3.745 214.955 3.995 215.965 ;
  LAYER M1 ;
        RECT 3.745 217.055 3.995 220.585 ;
  LAYER M1 ;
        RECT 3.745 220.835 3.995 221.845 ;
  LAYER M1 ;
        RECT 3.745 222.935 3.995 226.465 ;
  LAYER M1 ;
        RECT 3.745 226.715 3.995 227.725 ;
  LAYER M1 ;
        RECT 3.745 228.815 3.995 232.345 ;
  LAYER M1 ;
        RECT 3.745 232.595 3.995 233.605 ;
  LAYER M1 ;
        RECT 3.745 234.695 3.995 238.225 ;
  LAYER M1 ;
        RECT 3.745 238.475 3.995 239.485 ;
  LAYER M1 ;
        RECT 3.745 240.575 3.995 244.105 ;
  LAYER M1 ;
        RECT 3.745 244.355 3.995 245.365 ;
  LAYER M1 ;
        RECT 3.745 246.455 3.995 249.985 ;
  LAYER M1 ;
        RECT 3.745 250.235 3.995 251.245 ;
  LAYER M1 ;
        RECT 3.745 252.335 3.995 255.865 ;
  LAYER M1 ;
        RECT 3.745 256.115 3.995 257.125 ;
  LAYER M1 ;
        RECT 3.745 258.215 3.995 261.745 ;
  LAYER M1 ;
        RECT 3.745 261.995 3.995 263.005 ;
  LAYER M1 ;
        RECT 3.745 264.095 3.995 267.625 ;
  LAYER M1 ;
        RECT 3.745 267.875 3.995 268.885 ;
  LAYER M1 ;
        RECT 3.745 269.975 3.995 273.505 ;
  LAYER M1 ;
        RECT 3.745 273.755 3.995 274.765 ;
  LAYER M1 ;
        RECT 3.745 275.855 3.995 279.385 ;
  LAYER M1 ;
        RECT 3.745 279.635 3.995 280.645 ;
  LAYER M1 ;
        RECT 3.745 281.735 3.995 285.265 ;
  LAYER M1 ;
        RECT 3.745 285.515 3.995 286.525 ;
  LAYER M1 ;
        RECT 3.745 287.615 3.995 291.145 ;
  LAYER M1 ;
        RECT 3.745 291.395 3.995 292.405 ;
  LAYER M1 ;
        RECT 3.745 293.495 3.995 297.025 ;
  LAYER M1 ;
        RECT 3.745 297.275 3.995 298.285 ;
  LAYER M1 ;
        RECT 3.745 299.375 3.995 302.905 ;
  LAYER M1 ;
        RECT 3.745 303.155 3.995 304.165 ;
  LAYER M1 ;
        RECT 3.745 305.255 3.995 308.785 ;
  LAYER M1 ;
        RECT 3.745 309.035 3.995 310.045 ;
  LAYER M1 ;
        RECT 3.745 311.135 3.995 314.665 ;
  LAYER M1 ;
        RECT 3.745 314.915 3.995 315.925 ;
  LAYER M1 ;
        RECT 3.745 317.015 3.995 320.545 ;
  LAYER M1 ;
        RECT 3.745 320.795 3.995 321.805 ;
  LAYER M1 ;
        RECT 3.745 322.895 3.995 326.425 ;
  LAYER M1 ;
        RECT 3.745 326.675 3.995 327.685 ;
  LAYER M1 ;
        RECT 3.745 328.775 3.995 332.305 ;
  LAYER M1 ;
        RECT 3.745 332.555 3.995 333.565 ;
  LAYER M1 ;
        RECT 3.745 334.655 3.995 338.185 ;
  LAYER M1 ;
        RECT 3.745 338.435 3.995 339.445 ;
  LAYER M1 ;
        RECT 3.745 340.535 3.995 344.065 ;
  LAYER M1 ;
        RECT 3.745 344.315 3.995 345.325 ;
  LAYER M1 ;
        RECT 3.745 346.415 3.995 349.945 ;
  LAYER M1 ;
        RECT 3.745 350.195 3.995 351.205 ;
  LAYER M1 ;
        RECT 3.745 352.295 3.995 355.825 ;
  LAYER M1 ;
        RECT 3.745 356.075 3.995 357.085 ;
  LAYER M1 ;
        RECT 3.745 358.175 3.995 361.705 ;
  LAYER M1 ;
        RECT 3.745 361.955 3.995 362.965 ;
  LAYER M1 ;
        RECT 3.745 364.055 3.995 367.585 ;
  LAYER M1 ;
        RECT 3.745 367.835 3.995 368.845 ;
  LAYER M1 ;
        RECT 3.745 369.935 3.995 373.465 ;
  LAYER M1 ;
        RECT 3.745 373.715 3.995 374.725 ;
  LAYER M1 ;
        RECT 3.745 375.815 3.995 379.345 ;
  LAYER M1 ;
        RECT 3.745 379.595 3.995 380.605 ;
  LAYER M1 ;
        RECT 3.745 381.695 3.995 385.225 ;
  LAYER M1 ;
        RECT 3.745 385.475 3.995 386.485 ;
  LAYER M1 ;
        RECT 3.745 387.575 3.995 391.105 ;
  LAYER M1 ;
        RECT 3.745 391.355 3.995 392.365 ;
  LAYER M1 ;
        RECT 3.745 393.455 3.995 396.985 ;
  LAYER M1 ;
        RECT 3.745 397.235 3.995 398.245 ;
  LAYER M1 ;
        RECT 3.745 399.335 3.995 402.865 ;
  LAYER M1 ;
        RECT 3.745 403.115 3.995 404.125 ;
  LAYER M1 ;
        RECT 3.745 405.215 3.995 408.745 ;
  LAYER M1 ;
        RECT 3.745 408.995 3.995 410.005 ;
  LAYER M1 ;
        RECT 3.745 411.095 3.995 414.625 ;
  LAYER M1 ;
        RECT 3.745 414.875 3.995 415.885 ;
  LAYER M1 ;
        RECT 3.745 416.975 3.995 420.505 ;
  LAYER M1 ;
        RECT 3.745 420.755 3.995 421.765 ;
  LAYER M1 ;
        RECT 3.745 422.855 3.995 426.385 ;
  LAYER M1 ;
        RECT 3.745 426.635 3.995 427.645 ;
  LAYER M1 ;
        RECT 3.745 428.735 3.995 432.265 ;
  LAYER M1 ;
        RECT 3.745 432.515 3.995 433.525 ;
  LAYER M1 ;
        RECT 3.745 434.615 3.995 438.145 ;
  LAYER M1 ;
        RECT 3.745 438.395 3.995 439.405 ;
  LAYER M1 ;
        RECT 3.745 440.495 3.995 444.025 ;
  LAYER M1 ;
        RECT 3.745 444.275 3.995 445.285 ;
  LAYER M1 ;
        RECT 3.745 446.375 3.995 449.905 ;
  LAYER M1 ;
        RECT 3.745 450.155 3.995 451.165 ;
  LAYER M1 ;
        RECT 3.745 452.255 3.995 455.785 ;
  LAYER M1 ;
        RECT 3.745 456.035 3.995 457.045 ;
  LAYER M1 ;
        RECT 3.745 458.135 3.995 461.665 ;
  LAYER M1 ;
        RECT 3.745 461.915 3.995 462.925 ;
  LAYER M1 ;
        RECT 3.745 464.015 3.995 467.545 ;
  LAYER M1 ;
        RECT 3.745 467.795 3.995 468.805 ;
  LAYER M1 ;
        RECT 3.745 469.895 3.995 473.425 ;
  LAYER M1 ;
        RECT 3.745 473.675 3.995 474.685 ;
  LAYER M1 ;
        RECT 3.745 475.775 3.995 479.305 ;
  LAYER M1 ;
        RECT 3.745 479.555 3.995 480.565 ;
  LAYER M1 ;
        RECT 3.745 481.655 3.995 482.665 ;
  LAYER M1 ;
        RECT 3.315 64.175 3.565 67.705 ;
  LAYER M1 ;
        RECT 3.315 70.055 3.565 73.585 ;
  LAYER M1 ;
        RECT 3.315 75.935 3.565 79.465 ;
  LAYER M1 ;
        RECT 3.315 81.815 3.565 85.345 ;
  LAYER M1 ;
        RECT 3.315 87.695 3.565 91.225 ;
  LAYER M1 ;
        RECT 3.315 93.575 3.565 97.105 ;
  LAYER M1 ;
        RECT 3.315 99.455 3.565 102.985 ;
  LAYER M1 ;
        RECT 3.315 105.335 3.565 108.865 ;
  LAYER M1 ;
        RECT 3.315 111.215 3.565 114.745 ;
  LAYER M1 ;
        RECT 3.315 117.095 3.565 120.625 ;
  LAYER M1 ;
        RECT 3.315 122.975 3.565 126.505 ;
  LAYER M1 ;
        RECT 3.315 128.855 3.565 132.385 ;
  LAYER M1 ;
        RECT 3.315 134.735 3.565 138.265 ;
  LAYER M1 ;
        RECT 3.315 140.615 3.565 144.145 ;
  LAYER M1 ;
        RECT 3.315 146.495 3.565 150.025 ;
  LAYER M1 ;
        RECT 3.315 152.375 3.565 155.905 ;
  LAYER M1 ;
        RECT 3.315 158.255 3.565 161.785 ;
  LAYER M1 ;
        RECT 3.315 164.135 3.565 167.665 ;
  LAYER M1 ;
        RECT 3.315 170.015 3.565 173.545 ;
  LAYER M1 ;
        RECT 3.315 175.895 3.565 179.425 ;
  LAYER M1 ;
        RECT 3.315 181.775 3.565 185.305 ;
  LAYER M1 ;
        RECT 3.315 187.655 3.565 191.185 ;
  LAYER M1 ;
        RECT 3.315 193.535 3.565 197.065 ;
  LAYER M1 ;
        RECT 3.315 199.415 3.565 202.945 ;
  LAYER M1 ;
        RECT 3.315 205.295 3.565 208.825 ;
  LAYER M1 ;
        RECT 3.315 211.175 3.565 214.705 ;
  LAYER M1 ;
        RECT 3.315 217.055 3.565 220.585 ;
  LAYER M1 ;
        RECT 3.315 222.935 3.565 226.465 ;
  LAYER M1 ;
        RECT 3.315 228.815 3.565 232.345 ;
  LAYER M1 ;
        RECT 3.315 234.695 3.565 238.225 ;
  LAYER M1 ;
        RECT 3.315 240.575 3.565 244.105 ;
  LAYER M1 ;
        RECT 3.315 246.455 3.565 249.985 ;
  LAYER M1 ;
        RECT 3.315 252.335 3.565 255.865 ;
  LAYER M1 ;
        RECT 3.315 258.215 3.565 261.745 ;
  LAYER M1 ;
        RECT 3.315 264.095 3.565 267.625 ;
  LAYER M1 ;
        RECT 3.315 269.975 3.565 273.505 ;
  LAYER M1 ;
        RECT 3.315 275.855 3.565 279.385 ;
  LAYER M1 ;
        RECT 3.315 281.735 3.565 285.265 ;
  LAYER M1 ;
        RECT 3.315 287.615 3.565 291.145 ;
  LAYER M1 ;
        RECT 3.315 293.495 3.565 297.025 ;
  LAYER M1 ;
        RECT 3.315 299.375 3.565 302.905 ;
  LAYER M1 ;
        RECT 3.315 305.255 3.565 308.785 ;
  LAYER M1 ;
        RECT 3.315 311.135 3.565 314.665 ;
  LAYER M1 ;
        RECT 3.315 317.015 3.565 320.545 ;
  LAYER M1 ;
        RECT 3.315 322.895 3.565 326.425 ;
  LAYER M1 ;
        RECT 3.315 328.775 3.565 332.305 ;
  LAYER M1 ;
        RECT 3.315 334.655 3.565 338.185 ;
  LAYER M1 ;
        RECT 3.315 340.535 3.565 344.065 ;
  LAYER M1 ;
        RECT 3.315 346.415 3.565 349.945 ;
  LAYER M1 ;
        RECT 3.315 352.295 3.565 355.825 ;
  LAYER M1 ;
        RECT 3.315 358.175 3.565 361.705 ;
  LAYER M1 ;
        RECT 3.315 364.055 3.565 367.585 ;
  LAYER M1 ;
        RECT 3.315 369.935 3.565 373.465 ;
  LAYER M1 ;
        RECT 3.315 375.815 3.565 379.345 ;
  LAYER M1 ;
        RECT 3.315 381.695 3.565 385.225 ;
  LAYER M1 ;
        RECT 3.315 387.575 3.565 391.105 ;
  LAYER M1 ;
        RECT 3.315 393.455 3.565 396.985 ;
  LAYER M1 ;
        RECT 3.315 399.335 3.565 402.865 ;
  LAYER M1 ;
        RECT 3.315 405.215 3.565 408.745 ;
  LAYER M1 ;
        RECT 3.315 411.095 3.565 414.625 ;
  LAYER M1 ;
        RECT 3.315 416.975 3.565 420.505 ;
  LAYER M1 ;
        RECT 3.315 422.855 3.565 426.385 ;
  LAYER M1 ;
        RECT 3.315 428.735 3.565 432.265 ;
  LAYER M1 ;
        RECT 3.315 434.615 3.565 438.145 ;
  LAYER M1 ;
        RECT 3.315 440.495 3.565 444.025 ;
  LAYER M1 ;
        RECT 3.315 446.375 3.565 449.905 ;
  LAYER M1 ;
        RECT 3.315 452.255 3.565 455.785 ;
  LAYER M1 ;
        RECT 3.315 458.135 3.565 461.665 ;
  LAYER M1 ;
        RECT 3.315 464.015 3.565 467.545 ;
  LAYER M1 ;
        RECT 3.315 469.895 3.565 473.425 ;
  LAYER M1 ;
        RECT 3.315 475.775 3.565 479.305 ;
  LAYER M1 ;
        RECT 4.175 64.175 4.425 67.705 ;
  LAYER M1 ;
        RECT 4.175 70.055 4.425 73.585 ;
  LAYER M1 ;
        RECT 4.175 75.935 4.425 79.465 ;
  LAYER M1 ;
        RECT 4.175 81.815 4.425 85.345 ;
  LAYER M1 ;
        RECT 4.175 87.695 4.425 91.225 ;
  LAYER M1 ;
        RECT 4.175 93.575 4.425 97.105 ;
  LAYER M1 ;
        RECT 4.175 99.455 4.425 102.985 ;
  LAYER M1 ;
        RECT 4.175 105.335 4.425 108.865 ;
  LAYER M1 ;
        RECT 4.175 111.215 4.425 114.745 ;
  LAYER M1 ;
        RECT 4.175 117.095 4.425 120.625 ;
  LAYER M1 ;
        RECT 4.175 122.975 4.425 126.505 ;
  LAYER M1 ;
        RECT 4.175 128.855 4.425 132.385 ;
  LAYER M1 ;
        RECT 4.175 134.735 4.425 138.265 ;
  LAYER M1 ;
        RECT 4.175 140.615 4.425 144.145 ;
  LAYER M1 ;
        RECT 4.175 146.495 4.425 150.025 ;
  LAYER M1 ;
        RECT 4.175 152.375 4.425 155.905 ;
  LAYER M1 ;
        RECT 4.175 158.255 4.425 161.785 ;
  LAYER M1 ;
        RECT 4.175 164.135 4.425 167.665 ;
  LAYER M1 ;
        RECT 4.175 170.015 4.425 173.545 ;
  LAYER M1 ;
        RECT 4.175 175.895 4.425 179.425 ;
  LAYER M1 ;
        RECT 4.175 181.775 4.425 185.305 ;
  LAYER M1 ;
        RECT 4.175 187.655 4.425 191.185 ;
  LAYER M1 ;
        RECT 4.175 193.535 4.425 197.065 ;
  LAYER M1 ;
        RECT 4.175 199.415 4.425 202.945 ;
  LAYER M1 ;
        RECT 4.175 205.295 4.425 208.825 ;
  LAYER M1 ;
        RECT 4.175 211.175 4.425 214.705 ;
  LAYER M1 ;
        RECT 4.175 217.055 4.425 220.585 ;
  LAYER M1 ;
        RECT 4.175 222.935 4.425 226.465 ;
  LAYER M1 ;
        RECT 4.175 228.815 4.425 232.345 ;
  LAYER M1 ;
        RECT 4.175 234.695 4.425 238.225 ;
  LAYER M1 ;
        RECT 4.175 240.575 4.425 244.105 ;
  LAYER M1 ;
        RECT 4.175 246.455 4.425 249.985 ;
  LAYER M1 ;
        RECT 4.175 252.335 4.425 255.865 ;
  LAYER M1 ;
        RECT 4.175 258.215 4.425 261.745 ;
  LAYER M1 ;
        RECT 4.175 264.095 4.425 267.625 ;
  LAYER M1 ;
        RECT 4.175 269.975 4.425 273.505 ;
  LAYER M1 ;
        RECT 4.175 275.855 4.425 279.385 ;
  LAYER M1 ;
        RECT 4.175 281.735 4.425 285.265 ;
  LAYER M1 ;
        RECT 4.175 287.615 4.425 291.145 ;
  LAYER M1 ;
        RECT 4.175 293.495 4.425 297.025 ;
  LAYER M1 ;
        RECT 4.175 299.375 4.425 302.905 ;
  LAYER M1 ;
        RECT 4.175 305.255 4.425 308.785 ;
  LAYER M1 ;
        RECT 4.175 311.135 4.425 314.665 ;
  LAYER M1 ;
        RECT 4.175 317.015 4.425 320.545 ;
  LAYER M1 ;
        RECT 4.175 322.895 4.425 326.425 ;
  LAYER M1 ;
        RECT 4.175 328.775 4.425 332.305 ;
  LAYER M1 ;
        RECT 4.175 334.655 4.425 338.185 ;
  LAYER M1 ;
        RECT 4.175 340.535 4.425 344.065 ;
  LAYER M1 ;
        RECT 4.175 346.415 4.425 349.945 ;
  LAYER M1 ;
        RECT 4.175 352.295 4.425 355.825 ;
  LAYER M1 ;
        RECT 4.175 358.175 4.425 361.705 ;
  LAYER M1 ;
        RECT 4.175 364.055 4.425 367.585 ;
  LAYER M1 ;
        RECT 4.175 369.935 4.425 373.465 ;
  LAYER M1 ;
        RECT 4.175 375.815 4.425 379.345 ;
  LAYER M1 ;
        RECT 4.175 381.695 4.425 385.225 ;
  LAYER M1 ;
        RECT 4.175 387.575 4.425 391.105 ;
  LAYER M1 ;
        RECT 4.175 393.455 4.425 396.985 ;
  LAYER M1 ;
        RECT 4.175 399.335 4.425 402.865 ;
  LAYER M1 ;
        RECT 4.175 405.215 4.425 408.745 ;
  LAYER M1 ;
        RECT 4.175 411.095 4.425 414.625 ;
  LAYER M1 ;
        RECT 4.175 416.975 4.425 420.505 ;
  LAYER M1 ;
        RECT 4.175 422.855 4.425 426.385 ;
  LAYER M1 ;
        RECT 4.175 428.735 4.425 432.265 ;
  LAYER M1 ;
        RECT 4.175 434.615 4.425 438.145 ;
  LAYER M1 ;
        RECT 4.175 440.495 4.425 444.025 ;
  LAYER M1 ;
        RECT 4.175 446.375 4.425 449.905 ;
  LAYER M1 ;
        RECT 4.175 452.255 4.425 455.785 ;
  LAYER M1 ;
        RECT 4.175 458.135 4.425 461.665 ;
  LAYER M1 ;
        RECT 4.175 464.015 4.425 467.545 ;
  LAYER M1 ;
        RECT 4.175 469.895 4.425 473.425 ;
  LAYER M1 ;
        RECT 4.175 475.775 4.425 479.305 ;
  LAYER M2 ;
        RECT 2.84 64.12 4.04 64.4 ;
  LAYER M2 ;
        RECT 2.84 68.32 4.04 68.6 ;
  LAYER M2 ;
        RECT 3.27 64.54 4.47 64.82 ;
  LAYER M2 ;
        RECT 2.84 70 4.04 70.28 ;
  LAYER M2 ;
        RECT 2.84 74.2 4.04 74.48 ;
  LAYER M2 ;
        RECT 3.27 70.42 4.47 70.7 ;
  LAYER M2 ;
        RECT 2.84 75.88 4.04 76.16 ;
  LAYER M2 ;
        RECT 2.84 80.08 4.04 80.36 ;
  LAYER M2 ;
        RECT 3.27 76.3 4.47 76.58 ;
  LAYER M2 ;
        RECT 2.84 81.76 4.04 82.04 ;
  LAYER M2 ;
        RECT 2.84 85.96 4.04 86.24 ;
  LAYER M2 ;
        RECT 3.27 82.18 4.47 82.46 ;
  LAYER M2 ;
        RECT 2.84 87.64 4.04 87.92 ;
  LAYER M2 ;
        RECT 2.84 91.84 4.04 92.12 ;
  LAYER M2 ;
        RECT 3.27 88.06 4.47 88.34 ;
  LAYER M2 ;
        RECT 2.84 93.52 4.04 93.8 ;
  LAYER M2 ;
        RECT 2.84 97.72 4.04 98 ;
  LAYER M2 ;
        RECT 3.27 93.94 4.47 94.22 ;
  LAYER M2 ;
        RECT 2.84 99.4 4.04 99.68 ;
  LAYER M2 ;
        RECT 2.84 103.6 4.04 103.88 ;
  LAYER M2 ;
        RECT 3.27 99.82 4.47 100.1 ;
  LAYER M2 ;
        RECT 2.84 105.28 4.04 105.56 ;
  LAYER M2 ;
        RECT 2.84 109.48 4.04 109.76 ;
  LAYER M2 ;
        RECT 3.27 105.7 4.47 105.98 ;
  LAYER M2 ;
        RECT 2.84 111.16 4.04 111.44 ;
  LAYER M2 ;
        RECT 2.84 115.36 4.04 115.64 ;
  LAYER M2 ;
        RECT 3.27 111.58 4.47 111.86 ;
  LAYER M2 ;
        RECT 2.84 117.04 4.04 117.32 ;
  LAYER M2 ;
        RECT 2.84 121.24 4.04 121.52 ;
  LAYER M2 ;
        RECT 3.27 117.46 4.47 117.74 ;
  LAYER M2 ;
        RECT 2.84 122.92 4.04 123.2 ;
  LAYER M2 ;
        RECT 2.84 127.12 4.04 127.4 ;
  LAYER M2 ;
        RECT 3.27 123.34 4.47 123.62 ;
  LAYER M2 ;
        RECT 2.84 128.8 4.04 129.08 ;
  LAYER M2 ;
        RECT 2.84 133 4.04 133.28 ;
  LAYER M2 ;
        RECT 3.27 129.22 4.47 129.5 ;
  LAYER M2 ;
        RECT 2.84 134.68 4.04 134.96 ;
  LAYER M2 ;
        RECT 2.84 138.88 4.04 139.16 ;
  LAYER M2 ;
        RECT 3.27 135.1 4.47 135.38 ;
  LAYER M2 ;
        RECT 2.84 140.56 4.04 140.84 ;
  LAYER M2 ;
        RECT 2.84 144.76 4.04 145.04 ;
  LAYER M2 ;
        RECT 3.27 140.98 4.47 141.26 ;
  LAYER M2 ;
        RECT 2.84 146.44 4.04 146.72 ;
  LAYER M2 ;
        RECT 2.84 150.64 4.04 150.92 ;
  LAYER M2 ;
        RECT 3.27 146.86 4.47 147.14 ;
  LAYER M2 ;
        RECT 2.84 152.32 4.04 152.6 ;
  LAYER M2 ;
        RECT 2.84 156.52 4.04 156.8 ;
  LAYER M2 ;
        RECT 3.27 152.74 4.47 153.02 ;
  LAYER M2 ;
        RECT 2.84 158.2 4.04 158.48 ;
  LAYER M2 ;
        RECT 2.84 162.4 4.04 162.68 ;
  LAYER M2 ;
        RECT 3.27 158.62 4.47 158.9 ;
  LAYER M2 ;
        RECT 2.84 164.08 4.04 164.36 ;
  LAYER M2 ;
        RECT 2.84 168.28 4.04 168.56 ;
  LAYER M2 ;
        RECT 3.27 164.5 4.47 164.78 ;
  LAYER M2 ;
        RECT 2.84 169.96 4.04 170.24 ;
  LAYER M2 ;
        RECT 2.84 174.16 4.04 174.44 ;
  LAYER M2 ;
        RECT 3.27 170.38 4.47 170.66 ;
  LAYER M2 ;
        RECT 2.84 175.84 4.04 176.12 ;
  LAYER M2 ;
        RECT 2.84 180.04 4.04 180.32 ;
  LAYER M2 ;
        RECT 3.27 176.26 4.47 176.54 ;
  LAYER M2 ;
        RECT 2.84 181.72 4.04 182 ;
  LAYER M2 ;
        RECT 2.84 185.92 4.04 186.2 ;
  LAYER M2 ;
        RECT 3.27 182.14 4.47 182.42 ;
  LAYER M2 ;
        RECT 2.84 187.6 4.04 187.88 ;
  LAYER M2 ;
        RECT 2.84 191.8 4.04 192.08 ;
  LAYER M2 ;
        RECT 3.27 188.02 4.47 188.3 ;
  LAYER M2 ;
        RECT 2.84 193.48 4.04 193.76 ;
  LAYER M2 ;
        RECT 2.84 197.68 4.04 197.96 ;
  LAYER M2 ;
        RECT 3.27 193.9 4.47 194.18 ;
  LAYER M2 ;
        RECT 2.84 199.36 4.04 199.64 ;
  LAYER M2 ;
        RECT 2.84 203.56 4.04 203.84 ;
  LAYER M2 ;
        RECT 3.27 199.78 4.47 200.06 ;
  LAYER M2 ;
        RECT 2.84 205.24 4.04 205.52 ;
  LAYER M2 ;
        RECT 2.84 209.44 4.04 209.72 ;
  LAYER M2 ;
        RECT 3.27 205.66 4.47 205.94 ;
  LAYER M2 ;
        RECT 2.84 211.12 4.04 211.4 ;
  LAYER M2 ;
        RECT 2.84 215.32 4.04 215.6 ;
  LAYER M2 ;
        RECT 3.27 211.54 4.47 211.82 ;
  LAYER M2 ;
        RECT 2.84 217 4.04 217.28 ;
  LAYER M2 ;
        RECT 2.84 221.2 4.04 221.48 ;
  LAYER M2 ;
        RECT 3.27 217.42 4.47 217.7 ;
  LAYER M2 ;
        RECT 2.84 222.88 4.04 223.16 ;
  LAYER M2 ;
        RECT 2.84 227.08 4.04 227.36 ;
  LAYER M2 ;
        RECT 3.27 223.3 4.47 223.58 ;
  LAYER M2 ;
        RECT 2.84 228.76 4.04 229.04 ;
  LAYER M2 ;
        RECT 2.84 232.96 4.04 233.24 ;
  LAYER M2 ;
        RECT 3.27 229.18 4.47 229.46 ;
  LAYER M2 ;
        RECT 2.84 234.64 4.04 234.92 ;
  LAYER M2 ;
        RECT 2.84 238.84 4.04 239.12 ;
  LAYER M2 ;
        RECT 3.27 235.06 4.47 235.34 ;
  LAYER M2 ;
        RECT 2.84 240.52 4.04 240.8 ;
  LAYER M2 ;
        RECT 2.84 244.72 4.04 245 ;
  LAYER M2 ;
        RECT 3.27 240.94 4.47 241.22 ;
  LAYER M2 ;
        RECT 2.84 246.4 4.04 246.68 ;
  LAYER M2 ;
        RECT 2.84 250.6 4.04 250.88 ;
  LAYER M2 ;
        RECT 3.27 246.82 4.47 247.1 ;
  LAYER M2 ;
        RECT 2.84 252.28 4.04 252.56 ;
  LAYER M2 ;
        RECT 2.84 256.48 4.04 256.76 ;
  LAYER M2 ;
        RECT 3.27 252.7 4.47 252.98 ;
  LAYER M2 ;
        RECT 2.84 258.16 4.04 258.44 ;
  LAYER M2 ;
        RECT 2.84 262.36 4.04 262.64 ;
  LAYER M2 ;
        RECT 3.27 258.58 4.47 258.86 ;
  LAYER M2 ;
        RECT 2.84 264.04 4.04 264.32 ;
  LAYER M2 ;
        RECT 2.84 268.24 4.04 268.52 ;
  LAYER M2 ;
        RECT 3.27 264.46 4.47 264.74 ;
  LAYER M2 ;
        RECT 2.84 269.92 4.04 270.2 ;
  LAYER M2 ;
        RECT 2.84 274.12 4.04 274.4 ;
  LAYER M2 ;
        RECT 3.27 270.34 4.47 270.62 ;
  LAYER M2 ;
        RECT 2.84 275.8 4.04 276.08 ;
  LAYER M2 ;
        RECT 2.84 280 4.04 280.28 ;
  LAYER M2 ;
        RECT 3.27 276.22 4.47 276.5 ;
  LAYER M2 ;
        RECT 2.84 281.68 4.04 281.96 ;
  LAYER M2 ;
        RECT 2.84 285.88 4.04 286.16 ;
  LAYER M2 ;
        RECT 3.27 282.1 4.47 282.38 ;
  LAYER M2 ;
        RECT 2.84 287.56 4.04 287.84 ;
  LAYER M2 ;
        RECT 2.84 291.76 4.04 292.04 ;
  LAYER M2 ;
        RECT 3.27 287.98 4.47 288.26 ;
  LAYER M2 ;
        RECT 2.84 293.44 4.04 293.72 ;
  LAYER M2 ;
        RECT 2.84 297.64 4.04 297.92 ;
  LAYER M2 ;
        RECT 3.27 293.86 4.47 294.14 ;
  LAYER M2 ;
        RECT 2.84 299.32 4.04 299.6 ;
  LAYER M2 ;
        RECT 2.84 303.52 4.04 303.8 ;
  LAYER M2 ;
        RECT 3.27 299.74 4.47 300.02 ;
  LAYER M2 ;
        RECT 2.84 305.2 4.04 305.48 ;
  LAYER M2 ;
        RECT 2.84 309.4 4.04 309.68 ;
  LAYER M2 ;
        RECT 3.27 305.62 4.47 305.9 ;
  LAYER M2 ;
        RECT 2.84 311.08 4.04 311.36 ;
  LAYER M2 ;
        RECT 2.84 315.28 4.04 315.56 ;
  LAYER M2 ;
        RECT 3.27 311.5 4.47 311.78 ;
  LAYER M2 ;
        RECT 2.84 316.96 4.04 317.24 ;
  LAYER M2 ;
        RECT 2.84 321.16 4.04 321.44 ;
  LAYER M2 ;
        RECT 3.27 317.38 4.47 317.66 ;
  LAYER M2 ;
        RECT 2.84 322.84 4.04 323.12 ;
  LAYER M2 ;
        RECT 2.84 327.04 4.04 327.32 ;
  LAYER M2 ;
        RECT 3.27 323.26 4.47 323.54 ;
  LAYER M2 ;
        RECT 2.84 328.72 4.04 329 ;
  LAYER M2 ;
        RECT 2.84 332.92 4.04 333.2 ;
  LAYER M2 ;
        RECT 3.27 329.14 4.47 329.42 ;
  LAYER M2 ;
        RECT 2.84 334.6 4.04 334.88 ;
  LAYER M2 ;
        RECT 2.84 338.8 4.04 339.08 ;
  LAYER M2 ;
        RECT 3.27 335.02 4.47 335.3 ;
  LAYER M2 ;
        RECT 2.84 340.48 4.04 340.76 ;
  LAYER M2 ;
        RECT 2.84 344.68 4.04 344.96 ;
  LAYER M2 ;
        RECT 3.27 340.9 4.47 341.18 ;
  LAYER M2 ;
        RECT 2.84 346.36 4.04 346.64 ;
  LAYER M2 ;
        RECT 2.84 350.56 4.04 350.84 ;
  LAYER M2 ;
        RECT 3.27 346.78 4.47 347.06 ;
  LAYER M2 ;
        RECT 2.84 352.24 4.04 352.52 ;
  LAYER M2 ;
        RECT 2.84 356.44 4.04 356.72 ;
  LAYER M2 ;
        RECT 3.27 352.66 4.47 352.94 ;
  LAYER M2 ;
        RECT 2.84 358.12 4.04 358.4 ;
  LAYER M2 ;
        RECT 2.84 362.32 4.04 362.6 ;
  LAYER M2 ;
        RECT 3.27 358.54 4.47 358.82 ;
  LAYER M2 ;
        RECT 2.84 364 4.04 364.28 ;
  LAYER M2 ;
        RECT 2.84 368.2 4.04 368.48 ;
  LAYER M2 ;
        RECT 3.27 364.42 4.47 364.7 ;
  LAYER M2 ;
        RECT 2.84 369.88 4.04 370.16 ;
  LAYER M2 ;
        RECT 2.84 374.08 4.04 374.36 ;
  LAYER M2 ;
        RECT 3.27 370.3 4.47 370.58 ;
  LAYER M2 ;
        RECT 2.84 375.76 4.04 376.04 ;
  LAYER M2 ;
        RECT 2.84 379.96 4.04 380.24 ;
  LAYER M2 ;
        RECT 3.27 376.18 4.47 376.46 ;
  LAYER M2 ;
        RECT 2.84 381.64 4.04 381.92 ;
  LAYER M2 ;
        RECT 2.84 385.84 4.04 386.12 ;
  LAYER M2 ;
        RECT 3.27 382.06 4.47 382.34 ;
  LAYER M2 ;
        RECT 2.84 387.52 4.04 387.8 ;
  LAYER M2 ;
        RECT 2.84 391.72 4.04 392 ;
  LAYER M2 ;
        RECT 3.27 387.94 4.47 388.22 ;
  LAYER M2 ;
        RECT 2.84 393.4 4.04 393.68 ;
  LAYER M2 ;
        RECT 2.84 397.6 4.04 397.88 ;
  LAYER M2 ;
        RECT 3.27 393.82 4.47 394.1 ;
  LAYER M2 ;
        RECT 2.84 399.28 4.04 399.56 ;
  LAYER M2 ;
        RECT 2.84 403.48 4.04 403.76 ;
  LAYER M2 ;
        RECT 3.27 399.7 4.47 399.98 ;
  LAYER M2 ;
        RECT 2.84 405.16 4.04 405.44 ;
  LAYER M2 ;
        RECT 2.84 409.36 4.04 409.64 ;
  LAYER M2 ;
        RECT 3.27 405.58 4.47 405.86 ;
  LAYER M2 ;
        RECT 2.84 411.04 4.04 411.32 ;
  LAYER M2 ;
        RECT 2.84 415.24 4.04 415.52 ;
  LAYER M2 ;
        RECT 3.27 411.46 4.47 411.74 ;
  LAYER M2 ;
        RECT 2.84 416.92 4.04 417.2 ;
  LAYER M2 ;
        RECT 2.84 421.12 4.04 421.4 ;
  LAYER M2 ;
        RECT 3.27 417.34 4.47 417.62 ;
  LAYER M2 ;
        RECT 2.84 422.8 4.04 423.08 ;
  LAYER M2 ;
        RECT 2.84 427 4.04 427.28 ;
  LAYER M2 ;
        RECT 3.27 423.22 4.47 423.5 ;
  LAYER M2 ;
        RECT 2.84 428.68 4.04 428.96 ;
  LAYER M2 ;
        RECT 2.84 432.88 4.04 433.16 ;
  LAYER M2 ;
        RECT 3.27 429.1 4.47 429.38 ;
  LAYER M2 ;
        RECT 2.84 434.56 4.04 434.84 ;
  LAYER M2 ;
        RECT 2.84 438.76 4.04 439.04 ;
  LAYER M2 ;
        RECT 3.27 434.98 4.47 435.26 ;
  LAYER M2 ;
        RECT 2.84 440.44 4.04 440.72 ;
  LAYER M2 ;
        RECT 2.84 444.64 4.04 444.92 ;
  LAYER M2 ;
        RECT 3.27 440.86 4.47 441.14 ;
  LAYER M2 ;
        RECT 2.84 446.32 4.04 446.6 ;
  LAYER M2 ;
        RECT 2.84 450.52 4.04 450.8 ;
  LAYER M2 ;
        RECT 3.27 446.74 4.47 447.02 ;
  LAYER M2 ;
        RECT 2.84 452.2 4.04 452.48 ;
  LAYER M2 ;
        RECT 2.84 456.4 4.04 456.68 ;
  LAYER M2 ;
        RECT 3.27 452.62 4.47 452.9 ;
  LAYER M2 ;
        RECT 2.84 458.08 4.04 458.36 ;
  LAYER M2 ;
        RECT 2.84 462.28 4.04 462.56 ;
  LAYER M2 ;
        RECT 3.27 458.5 4.47 458.78 ;
  LAYER M2 ;
        RECT 2.84 463.96 4.04 464.24 ;
  LAYER M2 ;
        RECT 2.84 468.16 4.04 468.44 ;
  LAYER M2 ;
        RECT 3.27 464.38 4.47 464.66 ;
  LAYER M2 ;
        RECT 2.84 469.84 4.04 470.12 ;
  LAYER M2 ;
        RECT 2.84 474.04 4.04 474.32 ;
  LAYER M2 ;
        RECT 3.27 470.26 4.47 470.54 ;
  LAYER M2 ;
        RECT 2.84 475.72 4.04 476 ;
  LAYER M2 ;
        RECT 2.84 479.92 4.04 480.2 ;
  LAYER M2 ;
        RECT 3.27 476.14 4.47 476.42 ;
  LAYER M2 ;
        RECT 3.27 482.02 4.47 482.3 ;
  LAYER M3 ;
        RECT 3.73 64.1 4.01 480.22 ;
  LAYER M3 ;
        RECT 4.16 64.52 4.44 482.32 ;
  LAYER M1 ;
        RECT 1.165 56.615 1.415 60.145 ;
  LAYER M1 ;
        RECT 1.165 60.395 1.415 61.405 ;
  LAYER M1 ;
        RECT 1.165 62.495 1.415 63.505 ;
  LAYER M1 ;
        RECT 0.735 56.615 0.985 60.145 ;
  LAYER M1 ;
        RECT 1.595 56.615 1.845 60.145 ;
  LAYER M1 ;
        RECT 2.025 56.615 2.275 60.145 ;
  LAYER M1 ;
        RECT 2.025 60.395 2.275 61.405 ;
  LAYER M1 ;
        RECT 2.025 62.495 2.275 63.505 ;
  LAYER M1 ;
        RECT 2.455 56.615 2.705 60.145 ;
  LAYER M1 ;
        RECT 2.885 56.615 3.135 60.145 ;
  LAYER M1 ;
        RECT 2.885 60.395 3.135 61.405 ;
  LAYER M1 ;
        RECT 2.885 62.495 3.135 63.505 ;
  LAYER M1 ;
        RECT 3.315 56.615 3.565 60.145 ;
  LAYER M2 ;
        RECT 1.12 56.56 3.18 56.84 ;
  LAYER M2 ;
        RECT 1.12 60.76 3.18 61.04 ;
  LAYER M2 ;
        RECT 0.69 56.98 3.61 57.26 ;
  LAYER M2 ;
        RECT 1.12 62.86 3.18 63.14 ;
  LAYER M3 ;
        RECT 2.01 56.54 2.29 61.06 ;
  LAYER M3 ;
        RECT 2.44 56.96 2.72 63.16 ;
  LAYER M1 ;
        RECT 8.905 56.615 9.155 60.145 ;
  LAYER M1 ;
        RECT 8.905 60.395 9.155 61.405 ;
  LAYER M1 ;
        RECT 8.905 62.495 9.155 63.505 ;
  LAYER M1 ;
        RECT 9.335 56.615 9.585 60.145 ;
  LAYER M1 ;
        RECT 8.475 56.615 8.725 60.145 ;
  LAYER M1 ;
        RECT 8.045 56.615 8.295 60.145 ;
  LAYER M1 ;
        RECT 8.045 60.395 8.295 61.405 ;
  LAYER M1 ;
        RECT 8.045 62.495 8.295 63.505 ;
  LAYER M1 ;
        RECT 7.615 56.615 7.865 60.145 ;
  LAYER M1 ;
        RECT 7.185 56.615 7.435 60.145 ;
  LAYER M1 ;
        RECT 7.185 60.395 7.435 61.405 ;
  LAYER M1 ;
        RECT 7.185 62.495 7.435 63.505 ;
  LAYER M1 ;
        RECT 6.755 56.615 7.005 60.145 ;
  LAYER M2 ;
        RECT 7.14 56.56 9.2 56.84 ;
  LAYER M2 ;
        RECT 7.14 60.76 9.2 61.04 ;
  LAYER M2 ;
        RECT 6.71 56.98 9.63 57.26 ;
  LAYER M2 ;
        RECT 7.14 62.86 9.2 63.14 ;
  LAYER M3 ;
        RECT 8.03 56.54 8.31 61.06 ;
  LAYER M3 ;
        RECT 7.6 56.96 7.88 63.16 ;
  LAYER M1 ;
        RECT 6.325 64.175 6.575 67.705 ;
  LAYER M1 ;
        RECT 6.325 67.955 6.575 68.965 ;
  LAYER M1 ;
        RECT 6.325 70.055 6.575 73.585 ;
  LAYER M1 ;
        RECT 6.325 73.835 6.575 74.845 ;
  LAYER M1 ;
        RECT 6.325 75.935 6.575 79.465 ;
  LAYER M1 ;
        RECT 6.325 79.715 6.575 80.725 ;
  LAYER M1 ;
        RECT 6.325 81.815 6.575 85.345 ;
  LAYER M1 ;
        RECT 6.325 85.595 6.575 86.605 ;
  LAYER M1 ;
        RECT 6.325 87.695 6.575 91.225 ;
  LAYER M1 ;
        RECT 6.325 91.475 6.575 92.485 ;
  LAYER M1 ;
        RECT 6.325 93.575 6.575 97.105 ;
  LAYER M1 ;
        RECT 6.325 97.355 6.575 98.365 ;
  LAYER M1 ;
        RECT 6.325 99.455 6.575 102.985 ;
  LAYER M1 ;
        RECT 6.325 103.235 6.575 104.245 ;
  LAYER M1 ;
        RECT 6.325 105.335 6.575 108.865 ;
  LAYER M1 ;
        RECT 6.325 109.115 6.575 110.125 ;
  LAYER M1 ;
        RECT 6.325 111.215 6.575 114.745 ;
  LAYER M1 ;
        RECT 6.325 114.995 6.575 116.005 ;
  LAYER M1 ;
        RECT 6.325 117.095 6.575 120.625 ;
  LAYER M1 ;
        RECT 6.325 120.875 6.575 121.885 ;
  LAYER M1 ;
        RECT 6.325 122.975 6.575 126.505 ;
  LAYER M1 ;
        RECT 6.325 126.755 6.575 127.765 ;
  LAYER M1 ;
        RECT 6.325 128.855 6.575 132.385 ;
  LAYER M1 ;
        RECT 6.325 132.635 6.575 133.645 ;
  LAYER M1 ;
        RECT 6.325 134.735 6.575 138.265 ;
  LAYER M1 ;
        RECT 6.325 138.515 6.575 139.525 ;
  LAYER M1 ;
        RECT 6.325 140.615 6.575 144.145 ;
  LAYER M1 ;
        RECT 6.325 144.395 6.575 145.405 ;
  LAYER M1 ;
        RECT 6.325 146.495 6.575 150.025 ;
  LAYER M1 ;
        RECT 6.325 150.275 6.575 151.285 ;
  LAYER M1 ;
        RECT 6.325 152.375 6.575 155.905 ;
  LAYER M1 ;
        RECT 6.325 156.155 6.575 157.165 ;
  LAYER M1 ;
        RECT 6.325 158.255 6.575 161.785 ;
  LAYER M1 ;
        RECT 6.325 162.035 6.575 163.045 ;
  LAYER M1 ;
        RECT 6.325 164.135 6.575 167.665 ;
  LAYER M1 ;
        RECT 6.325 167.915 6.575 168.925 ;
  LAYER M1 ;
        RECT 6.325 170.015 6.575 173.545 ;
  LAYER M1 ;
        RECT 6.325 173.795 6.575 174.805 ;
  LAYER M1 ;
        RECT 6.325 175.895 6.575 179.425 ;
  LAYER M1 ;
        RECT 6.325 179.675 6.575 180.685 ;
  LAYER M1 ;
        RECT 6.325 181.775 6.575 185.305 ;
  LAYER M1 ;
        RECT 6.325 185.555 6.575 186.565 ;
  LAYER M1 ;
        RECT 6.325 187.655 6.575 191.185 ;
  LAYER M1 ;
        RECT 6.325 191.435 6.575 192.445 ;
  LAYER M1 ;
        RECT 6.325 193.535 6.575 197.065 ;
  LAYER M1 ;
        RECT 6.325 197.315 6.575 198.325 ;
  LAYER M1 ;
        RECT 6.325 199.415 6.575 202.945 ;
  LAYER M1 ;
        RECT 6.325 203.195 6.575 204.205 ;
  LAYER M1 ;
        RECT 6.325 205.295 6.575 208.825 ;
  LAYER M1 ;
        RECT 6.325 209.075 6.575 210.085 ;
  LAYER M1 ;
        RECT 6.325 211.175 6.575 214.705 ;
  LAYER M1 ;
        RECT 6.325 214.955 6.575 215.965 ;
  LAYER M1 ;
        RECT 6.325 217.055 6.575 220.585 ;
  LAYER M1 ;
        RECT 6.325 220.835 6.575 221.845 ;
  LAYER M1 ;
        RECT 6.325 222.935 6.575 226.465 ;
  LAYER M1 ;
        RECT 6.325 226.715 6.575 227.725 ;
  LAYER M1 ;
        RECT 6.325 228.815 6.575 232.345 ;
  LAYER M1 ;
        RECT 6.325 232.595 6.575 233.605 ;
  LAYER M1 ;
        RECT 6.325 234.695 6.575 238.225 ;
  LAYER M1 ;
        RECT 6.325 238.475 6.575 239.485 ;
  LAYER M1 ;
        RECT 6.325 240.575 6.575 244.105 ;
  LAYER M1 ;
        RECT 6.325 244.355 6.575 245.365 ;
  LAYER M1 ;
        RECT 6.325 246.455 6.575 249.985 ;
  LAYER M1 ;
        RECT 6.325 250.235 6.575 251.245 ;
  LAYER M1 ;
        RECT 6.325 252.335 6.575 255.865 ;
  LAYER M1 ;
        RECT 6.325 256.115 6.575 257.125 ;
  LAYER M1 ;
        RECT 6.325 258.215 6.575 261.745 ;
  LAYER M1 ;
        RECT 6.325 261.995 6.575 263.005 ;
  LAYER M1 ;
        RECT 6.325 264.095 6.575 267.625 ;
  LAYER M1 ;
        RECT 6.325 267.875 6.575 268.885 ;
  LAYER M1 ;
        RECT 6.325 269.975 6.575 273.505 ;
  LAYER M1 ;
        RECT 6.325 273.755 6.575 274.765 ;
  LAYER M1 ;
        RECT 6.325 275.855 6.575 279.385 ;
  LAYER M1 ;
        RECT 6.325 279.635 6.575 280.645 ;
  LAYER M1 ;
        RECT 6.325 281.735 6.575 285.265 ;
  LAYER M1 ;
        RECT 6.325 285.515 6.575 286.525 ;
  LAYER M1 ;
        RECT 6.325 287.615 6.575 291.145 ;
  LAYER M1 ;
        RECT 6.325 291.395 6.575 292.405 ;
  LAYER M1 ;
        RECT 6.325 293.495 6.575 297.025 ;
  LAYER M1 ;
        RECT 6.325 297.275 6.575 298.285 ;
  LAYER M1 ;
        RECT 6.325 299.375 6.575 302.905 ;
  LAYER M1 ;
        RECT 6.325 303.155 6.575 304.165 ;
  LAYER M1 ;
        RECT 6.325 305.255 6.575 308.785 ;
  LAYER M1 ;
        RECT 6.325 309.035 6.575 310.045 ;
  LAYER M1 ;
        RECT 6.325 311.135 6.575 314.665 ;
  LAYER M1 ;
        RECT 6.325 314.915 6.575 315.925 ;
  LAYER M1 ;
        RECT 6.325 317.015 6.575 320.545 ;
  LAYER M1 ;
        RECT 6.325 320.795 6.575 321.805 ;
  LAYER M1 ;
        RECT 6.325 322.895 6.575 326.425 ;
  LAYER M1 ;
        RECT 6.325 326.675 6.575 327.685 ;
  LAYER M1 ;
        RECT 6.325 328.775 6.575 332.305 ;
  LAYER M1 ;
        RECT 6.325 332.555 6.575 333.565 ;
  LAYER M1 ;
        RECT 6.325 334.655 6.575 338.185 ;
  LAYER M1 ;
        RECT 6.325 338.435 6.575 339.445 ;
  LAYER M1 ;
        RECT 6.325 340.535 6.575 344.065 ;
  LAYER M1 ;
        RECT 6.325 344.315 6.575 345.325 ;
  LAYER M1 ;
        RECT 6.325 346.415 6.575 349.945 ;
  LAYER M1 ;
        RECT 6.325 350.195 6.575 351.205 ;
  LAYER M1 ;
        RECT 6.325 352.295 6.575 355.825 ;
  LAYER M1 ;
        RECT 6.325 356.075 6.575 357.085 ;
  LAYER M1 ;
        RECT 6.325 358.175 6.575 361.705 ;
  LAYER M1 ;
        RECT 6.325 361.955 6.575 362.965 ;
  LAYER M1 ;
        RECT 6.325 364.055 6.575 367.585 ;
  LAYER M1 ;
        RECT 6.325 367.835 6.575 368.845 ;
  LAYER M1 ;
        RECT 6.325 369.935 6.575 373.465 ;
  LAYER M1 ;
        RECT 6.325 373.715 6.575 374.725 ;
  LAYER M1 ;
        RECT 6.325 375.815 6.575 379.345 ;
  LAYER M1 ;
        RECT 6.325 379.595 6.575 380.605 ;
  LAYER M1 ;
        RECT 6.325 381.695 6.575 385.225 ;
  LAYER M1 ;
        RECT 6.325 385.475 6.575 386.485 ;
  LAYER M1 ;
        RECT 6.325 387.575 6.575 391.105 ;
  LAYER M1 ;
        RECT 6.325 391.355 6.575 392.365 ;
  LAYER M1 ;
        RECT 6.325 393.455 6.575 396.985 ;
  LAYER M1 ;
        RECT 6.325 397.235 6.575 398.245 ;
  LAYER M1 ;
        RECT 6.325 399.335 6.575 402.865 ;
  LAYER M1 ;
        RECT 6.325 403.115 6.575 404.125 ;
  LAYER M1 ;
        RECT 6.325 405.215 6.575 408.745 ;
  LAYER M1 ;
        RECT 6.325 408.995 6.575 410.005 ;
  LAYER M1 ;
        RECT 6.325 411.095 6.575 414.625 ;
  LAYER M1 ;
        RECT 6.325 414.875 6.575 415.885 ;
  LAYER M1 ;
        RECT 6.325 416.975 6.575 420.505 ;
  LAYER M1 ;
        RECT 6.325 420.755 6.575 421.765 ;
  LAYER M1 ;
        RECT 6.325 422.855 6.575 426.385 ;
  LAYER M1 ;
        RECT 6.325 426.635 6.575 427.645 ;
  LAYER M1 ;
        RECT 6.325 428.735 6.575 432.265 ;
  LAYER M1 ;
        RECT 6.325 432.515 6.575 433.525 ;
  LAYER M1 ;
        RECT 6.325 434.615 6.575 438.145 ;
  LAYER M1 ;
        RECT 6.325 438.395 6.575 439.405 ;
  LAYER M1 ;
        RECT 6.325 440.495 6.575 444.025 ;
  LAYER M1 ;
        RECT 6.325 444.275 6.575 445.285 ;
  LAYER M1 ;
        RECT 6.325 446.375 6.575 449.905 ;
  LAYER M1 ;
        RECT 6.325 450.155 6.575 451.165 ;
  LAYER M1 ;
        RECT 6.325 452.255 6.575 455.785 ;
  LAYER M1 ;
        RECT 6.325 456.035 6.575 457.045 ;
  LAYER M1 ;
        RECT 6.325 458.135 6.575 461.665 ;
  LAYER M1 ;
        RECT 6.325 461.915 6.575 462.925 ;
  LAYER M1 ;
        RECT 6.325 464.015 6.575 467.545 ;
  LAYER M1 ;
        RECT 6.325 467.795 6.575 468.805 ;
  LAYER M1 ;
        RECT 6.325 469.895 6.575 473.425 ;
  LAYER M1 ;
        RECT 6.325 473.675 6.575 474.685 ;
  LAYER M1 ;
        RECT 6.325 475.775 6.575 479.305 ;
  LAYER M1 ;
        RECT 6.325 479.555 6.575 480.565 ;
  LAYER M1 ;
        RECT 6.325 481.655 6.575 482.665 ;
  LAYER M1 ;
        RECT 6.755 64.175 7.005 67.705 ;
  LAYER M1 ;
        RECT 6.755 70.055 7.005 73.585 ;
  LAYER M1 ;
        RECT 6.755 75.935 7.005 79.465 ;
  LAYER M1 ;
        RECT 6.755 81.815 7.005 85.345 ;
  LAYER M1 ;
        RECT 6.755 87.695 7.005 91.225 ;
  LAYER M1 ;
        RECT 6.755 93.575 7.005 97.105 ;
  LAYER M1 ;
        RECT 6.755 99.455 7.005 102.985 ;
  LAYER M1 ;
        RECT 6.755 105.335 7.005 108.865 ;
  LAYER M1 ;
        RECT 6.755 111.215 7.005 114.745 ;
  LAYER M1 ;
        RECT 6.755 117.095 7.005 120.625 ;
  LAYER M1 ;
        RECT 6.755 122.975 7.005 126.505 ;
  LAYER M1 ;
        RECT 6.755 128.855 7.005 132.385 ;
  LAYER M1 ;
        RECT 6.755 134.735 7.005 138.265 ;
  LAYER M1 ;
        RECT 6.755 140.615 7.005 144.145 ;
  LAYER M1 ;
        RECT 6.755 146.495 7.005 150.025 ;
  LAYER M1 ;
        RECT 6.755 152.375 7.005 155.905 ;
  LAYER M1 ;
        RECT 6.755 158.255 7.005 161.785 ;
  LAYER M1 ;
        RECT 6.755 164.135 7.005 167.665 ;
  LAYER M1 ;
        RECT 6.755 170.015 7.005 173.545 ;
  LAYER M1 ;
        RECT 6.755 175.895 7.005 179.425 ;
  LAYER M1 ;
        RECT 6.755 181.775 7.005 185.305 ;
  LAYER M1 ;
        RECT 6.755 187.655 7.005 191.185 ;
  LAYER M1 ;
        RECT 6.755 193.535 7.005 197.065 ;
  LAYER M1 ;
        RECT 6.755 199.415 7.005 202.945 ;
  LAYER M1 ;
        RECT 6.755 205.295 7.005 208.825 ;
  LAYER M1 ;
        RECT 6.755 211.175 7.005 214.705 ;
  LAYER M1 ;
        RECT 6.755 217.055 7.005 220.585 ;
  LAYER M1 ;
        RECT 6.755 222.935 7.005 226.465 ;
  LAYER M1 ;
        RECT 6.755 228.815 7.005 232.345 ;
  LAYER M1 ;
        RECT 6.755 234.695 7.005 238.225 ;
  LAYER M1 ;
        RECT 6.755 240.575 7.005 244.105 ;
  LAYER M1 ;
        RECT 6.755 246.455 7.005 249.985 ;
  LAYER M1 ;
        RECT 6.755 252.335 7.005 255.865 ;
  LAYER M1 ;
        RECT 6.755 258.215 7.005 261.745 ;
  LAYER M1 ;
        RECT 6.755 264.095 7.005 267.625 ;
  LAYER M1 ;
        RECT 6.755 269.975 7.005 273.505 ;
  LAYER M1 ;
        RECT 6.755 275.855 7.005 279.385 ;
  LAYER M1 ;
        RECT 6.755 281.735 7.005 285.265 ;
  LAYER M1 ;
        RECT 6.755 287.615 7.005 291.145 ;
  LAYER M1 ;
        RECT 6.755 293.495 7.005 297.025 ;
  LAYER M1 ;
        RECT 6.755 299.375 7.005 302.905 ;
  LAYER M1 ;
        RECT 6.755 305.255 7.005 308.785 ;
  LAYER M1 ;
        RECT 6.755 311.135 7.005 314.665 ;
  LAYER M1 ;
        RECT 6.755 317.015 7.005 320.545 ;
  LAYER M1 ;
        RECT 6.755 322.895 7.005 326.425 ;
  LAYER M1 ;
        RECT 6.755 328.775 7.005 332.305 ;
  LAYER M1 ;
        RECT 6.755 334.655 7.005 338.185 ;
  LAYER M1 ;
        RECT 6.755 340.535 7.005 344.065 ;
  LAYER M1 ;
        RECT 6.755 346.415 7.005 349.945 ;
  LAYER M1 ;
        RECT 6.755 352.295 7.005 355.825 ;
  LAYER M1 ;
        RECT 6.755 358.175 7.005 361.705 ;
  LAYER M1 ;
        RECT 6.755 364.055 7.005 367.585 ;
  LAYER M1 ;
        RECT 6.755 369.935 7.005 373.465 ;
  LAYER M1 ;
        RECT 6.755 375.815 7.005 379.345 ;
  LAYER M1 ;
        RECT 6.755 381.695 7.005 385.225 ;
  LAYER M1 ;
        RECT 6.755 387.575 7.005 391.105 ;
  LAYER M1 ;
        RECT 6.755 393.455 7.005 396.985 ;
  LAYER M1 ;
        RECT 6.755 399.335 7.005 402.865 ;
  LAYER M1 ;
        RECT 6.755 405.215 7.005 408.745 ;
  LAYER M1 ;
        RECT 6.755 411.095 7.005 414.625 ;
  LAYER M1 ;
        RECT 6.755 416.975 7.005 420.505 ;
  LAYER M1 ;
        RECT 6.755 422.855 7.005 426.385 ;
  LAYER M1 ;
        RECT 6.755 428.735 7.005 432.265 ;
  LAYER M1 ;
        RECT 6.755 434.615 7.005 438.145 ;
  LAYER M1 ;
        RECT 6.755 440.495 7.005 444.025 ;
  LAYER M1 ;
        RECT 6.755 446.375 7.005 449.905 ;
  LAYER M1 ;
        RECT 6.755 452.255 7.005 455.785 ;
  LAYER M1 ;
        RECT 6.755 458.135 7.005 461.665 ;
  LAYER M1 ;
        RECT 6.755 464.015 7.005 467.545 ;
  LAYER M1 ;
        RECT 6.755 469.895 7.005 473.425 ;
  LAYER M1 ;
        RECT 6.755 475.775 7.005 479.305 ;
  LAYER M1 ;
        RECT 5.895 64.175 6.145 67.705 ;
  LAYER M1 ;
        RECT 5.895 70.055 6.145 73.585 ;
  LAYER M1 ;
        RECT 5.895 75.935 6.145 79.465 ;
  LAYER M1 ;
        RECT 5.895 81.815 6.145 85.345 ;
  LAYER M1 ;
        RECT 5.895 87.695 6.145 91.225 ;
  LAYER M1 ;
        RECT 5.895 93.575 6.145 97.105 ;
  LAYER M1 ;
        RECT 5.895 99.455 6.145 102.985 ;
  LAYER M1 ;
        RECT 5.895 105.335 6.145 108.865 ;
  LAYER M1 ;
        RECT 5.895 111.215 6.145 114.745 ;
  LAYER M1 ;
        RECT 5.895 117.095 6.145 120.625 ;
  LAYER M1 ;
        RECT 5.895 122.975 6.145 126.505 ;
  LAYER M1 ;
        RECT 5.895 128.855 6.145 132.385 ;
  LAYER M1 ;
        RECT 5.895 134.735 6.145 138.265 ;
  LAYER M1 ;
        RECT 5.895 140.615 6.145 144.145 ;
  LAYER M1 ;
        RECT 5.895 146.495 6.145 150.025 ;
  LAYER M1 ;
        RECT 5.895 152.375 6.145 155.905 ;
  LAYER M1 ;
        RECT 5.895 158.255 6.145 161.785 ;
  LAYER M1 ;
        RECT 5.895 164.135 6.145 167.665 ;
  LAYER M1 ;
        RECT 5.895 170.015 6.145 173.545 ;
  LAYER M1 ;
        RECT 5.895 175.895 6.145 179.425 ;
  LAYER M1 ;
        RECT 5.895 181.775 6.145 185.305 ;
  LAYER M1 ;
        RECT 5.895 187.655 6.145 191.185 ;
  LAYER M1 ;
        RECT 5.895 193.535 6.145 197.065 ;
  LAYER M1 ;
        RECT 5.895 199.415 6.145 202.945 ;
  LAYER M1 ;
        RECT 5.895 205.295 6.145 208.825 ;
  LAYER M1 ;
        RECT 5.895 211.175 6.145 214.705 ;
  LAYER M1 ;
        RECT 5.895 217.055 6.145 220.585 ;
  LAYER M1 ;
        RECT 5.895 222.935 6.145 226.465 ;
  LAYER M1 ;
        RECT 5.895 228.815 6.145 232.345 ;
  LAYER M1 ;
        RECT 5.895 234.695 6.145 238.225 ;
  LAYER M1 ;
        RECT 5.895 240.575 6.145 244.105 ;
  LAYER M1 ;
        RECT 5.895 246.455 6.145 249.985 ;
  LAYER M1 ;
        RECT 5.895 252.335 6.145 255.865 ;
  LAYER M1 ;
        RECT 5.895 258.215 6.145 261.745 ;
  LAYER M1 ;
        RECT 5.895 264.095 6.145 267.625 ;
  LAYER M1 ;
        RECT 5.895 269.975 6.145 273.505 ;
  LAYER M1 ;
        RECT 5.895 275.855 6.145 279.385 ;
  LAYER M1 ;
        RECT 5.895 281.735 6.145 285.265 ;
  LAYER M1 ;
        RECT 5.895 287.615 6.145 291.145 ;
  LAYER M1 ;
        RECT 5.895 293.495 6.145 297.025 ;
  LAYER M1 ;
        RECT 5.895 299.375 6.145 302.905 ;
  LAYER M1 ;
        RECT 5.895 305.255 6.145 308.785 ;
  LAYER M1 ;
        RECT 5.895 311.135 6.145 314.665 ;
  LAYER M1 ;
        RECT 5.895 317.015 6.145 320.545 ;
  LAYER M1 ;
        RECT 5.895 322.895 6.145 326.425 ;
  LAYER M1 ;
        RECT 5.895 328.775 6.145 332.305 ;
  LAYER M1 ;
        RECT 5.895 334.655 6.145 338.185 ;
  LAYER M1 ;
        RECT 5.895 340.535 6.145 344.065 ;
  LAYER M1 ;
        RECT 5.895 346.415 6.145 349.945 ;
  LAYER M1 ;
        RECT 5.895 352.295 6.145 355.825 ;
  LAYER M1 ;
        RECT 5.895 358.175 6.145 361.705 ;
  LAYER M1 ;
        RECT 5.895 364.055 6.145 367.585 ;
  LAYER M1 ;
        RECT 5.895 369.935 6.145 373.465 ;
  LAYER M1 ;
        RECT 5.895 375.815 6.145 379.345 ;
  LAYER M1 ;
        RECT 5.895 381.695 6.145 385.225 ;
  LAYER M1 ;
        RECT 5.895 387.575 6.145 391.105 ;
  LAYER M1 ;
        RECT 5.895 393.455 6.145 396.985 ;
  LAYER M1 ;
        RECT 5.895 399.335 6.145 402.865 ;
  LAYER M1 ;
        RECT 5.895 405.215 6.145 408.745 ;
  LAYER M1 ;
        RECT 5.895 411.095 6.145 414.625 ;
  LAYER M1 ;
        RECT 5.895 416.975 6.145 420.505 ;
  LAYER M1 ;
        RECT 5.895 422.855 6.145 426.385 ;
  LAYER M1 ;
        RECT 5.895 428.735 6.145 432.265 ;
  LAYER M1 ;
        RECT 5.895 434.615 6.145 438.145 ;
  LAYER M1 ;
        RECT 5.895 440.495 6.145 444.025 ;
  LAYER M1 ;
        RECT 5.895 446.375 6.145 449.905 ;
  LAYER M1 ;
        RECT 5.895 452.255 6.145 455.785 ;
  LAYER M1 ;
        RECT 5.895 458.135 6.145 461.665 ;
  LAYER M1 ;
        RECT 5.895 464.015 6.145 467.545 ;
  LAYER M1 ;
        RECT 5.895 469.895 6.145 473.425 ;
  LAYER M1 ;
        RECT 5.895 475.775 6.145 479.305 ;
  LAYER M2 ;
        RECT 6.28 64.12 7.48 64.4 ;
  LAYER M2 ;
        RECT 6.28 68.32 7.48 68.6 ;
  LAYER M2 ;
        RECT 5.85 64.54 7.05 64.82 ;
  LAYER M2 ;
        RECT 6.28 70 7.48 70.28 ;
  LAYER M2 ;
        RECT 6.28 74.2 7.48 74.48 ;
  LAYER M2 ;
        RECT 5.85 70.42 7.05 70.7 ;
  LAYER M2 ;
        RECT 6.28 75.88 7.48 76.16 ;
  LAYER M2 ;
        RECT 6.28 80.08 7.48 80.36 ;
  LAYER M2 ;
        RECT 5.85 76.3 7.05 76.58 ;
  LAYER M2 ;
        RECT 6.28 81.76 7.48 82.04 ;
  LAYER M2 ;
        RECT 6.28 85.96 7.48 86.24 ;
  LAYER M2 ;
        RECT 5.85 82.18 7.05 82.46 ;
  LAYER M2 ;
        RECT 6.28 87.64 7.48 87.92 ;
  LAYER M2 ;
        RECT 6.28 91.84 7.48 92.12 ;
  LAYER M2 ;
        RECT 5.85 88.06 7.05 88.34 ;
  LAYER M2 ;
        RECT 6.28 93.52 7.48 93.8 ;
  LAYER M2 ;
        RECT 6.28 97.72 7.48 98 ;
  LAYER M2 ;
        RECT 5.85 93.94 7.05 94.22 ;
  LAYER M2 ;
        RECT 6.28 99.4 7.48 99.68 ;
  LAYER M2 ;
        RECT 6.28 103.6 7.48 103.88 ;
  LAYER M2 ;
        RECT 5.85 99.82 7.05 100.1 ;
  LAYER M2 ;
        RECT 6.28 105.28 7.48 105.56 ;
  LAYER M2 ;
        RECT 6.28 109.48 7.48 109.76 ;
  LAYER M2 ;
        RECT 5.85 105.7 7.05 105.98 ;
  LAYER M2 ;
        RECT 6.28 111.16 7.48 111.44 ;
  LAYER M2 ;
        RECT 6.28 115.36 7.48 115.64 ;
  LAYER M2 ;
        RECT 5.85 111.58 7.05 111.86 ;
  LAYER M2 ;
        RECT 6.28 117.04 7.48 117.32 ;
  LAYER M2 ;
        RECT 6.28 121.24 7.48 121.52 ;
  LAYER M2 ;
        RECT 5.85 117.46 7.05 117.74 ;
  LAYER M2 ;
        RECT 6.28 122.92 7.48 123.2 ;
  LAYER M2 ;
        RECT 6.28 127.12 7.48 127.4 ;
  LAYER M2 ;
        RECT 5.85 123.34 7.05 123.62 ;
  LAYER M2 ;
        RECT 6.28 128.8 7.48 129.08 ;
  LAYER M2 ;
        RECT 6.28 133 7.48 133.28 ;
  LAYER M2 ;
        RECT 5.85 129.22 7.05 129.5 ;
  LAYER M2 ;
        RECT 6.28 134.68 7.48 134.96 ;
  LAYER M2 ;
        RECT 6.28 138.88 7.48 139.16 ;
  LAYER M2 ;
        RECT 5.85 135.1 7.05 135.38 ;
  LAYER M2 ;
        RECT 6.28 140.56 7.48 140.84 ;
  LAYER M2 ;
        RECT 6.28 144.76 7.48 145.04 ;
  LAYER M2 ;
        RECT 5.85 140.98 7.05 141.26 ;
  LAYER M2 ;
        RECT 6.28 146.44 7.48 146.72 ;
  LAYER M2 ;
        RECT 6.28 150.64 7.48 150.92 ;
  LAYER M2 ;
        RECT 5.85 146.86 7.05 147.14 ;
  LAYER M2 ;
        RECT 6.28 152.32 7.48 152.6 ;
  LAYER M2 ;
        RECT 6.28 156.52 7.48 156.8 ;
  LAYER M2 ;
        RECT 5.85 152.74 7.05 153.02 ;
  LAYER M2 ;
        RECT 6.28 158.2 7.48 158.48 ;
  LAYER M2 ;
        RECT 6.28 162.4 7.48 162.68 ;
  LAYER M2 ;
        RECT 5.85 158.62 7.05 158.9 ;
  LAYER M2 ;
        RECT 6.28 164.08 7.48 164.36 ;
  LAYER M2 ;
        RECT 6.28 168.28 7.48 168.56 ;
  LAYER M2 ;
        RECT 5.85 164.5 7.05 164.78 ;
  LAYER M2 ;
        RECT 6.28 169.96 7.48 170.24 ;
  LAYER M2 ;
        RECT 6.28 174.16 7.48 174.44 ;
  LAYER M2 ;
        RECT 5.85 170.38 7.05 170.66 ;
  LAYER M2 ;
        RECT 6.28 175.84 7.48 176.12 ;
  LAYER M2 ;
        RECT 6.28 180.04 7.48 180.32 ;
  LAYER M2 ;
        RECT 5.85 176.26 7.05 176.54 ;
  LAYER M2 ;
        RECT 6.28 181.72 7.48 182 ;
  LAYER M2 ;
        RECT 6.28 185.92 7.48 186.2 ;
  LAYER M2 ;
        RECT 5.85 182.14 7.05 182.42 ;
  LAYER M2 ;
        RECT 6.28 187.6 7.48 187.88 ;
  LAYER M2 ;
        RECT 6.28 191.8 7.48 192.08 ;
  LAYER M2 ;
        RECT 5.85 188.02 7.05 188.3 ;
  LAYER M2 ;
        RECT 6.28 193.48 7.48 193.76 ;
  LAYER M2 ;
        RECT 6.28 197.68 7.48 197.96 ;
  LAYER M2 ;
        RECT 5.85 193.9 7.05 194.18 ;
  LAYER M2 ;
        RECT 6.28 199.36 7.48 199.64 ;
  LAYER M2 ;
        RECT 6.28 203.56 7.48 203.84 ;
  LAYER M2 ;
        RECT 5.85 199.78 7.05 200.06 ;
  LAYER M2 ;
        RECT 6.28 205.24 7.48 205.52 ;
  LAYER M2 ;
        RECT 6.28 209.44 7.48 209.72 ;
  LAYER M2 ;
        RECT 5.85 205.66 7.05 205.94 ;
  LAYER M2 ;
        RECT 6.28 211.12 7.48 211.4 ;
  LAYER M2 ;
        RECT 6.28 215.32 7.48 215.6 ;
  LAYER M2 ;
        RECT 5.85 211.54 7.05 211.82 ;
  LAYER M2 ;
        RECT 6.28 217 7.48 217.28 ;
  LAYER M2 ;
        RECT 6.28 221.2 7.48 221.48 ;
  LAYER M2 ;
        RECT 5.85 217.42 7.05 217.7 ;
  LAYER M2 ;
        RECT 6.28 222.88 7.48 223.16 ;
  LAYER M2 ;
        RECT 6.28 227.08 7.48 227.36 ;
  LAYER M2 ;
        RECT 5.85 223.3 7.05 223.58 ;
  LAYER M2 ;
        RECT 6.28 228.76 7.48 229.04 ;
  LAYER M2 ;
        RECT 6.28 232.96 7.48 233.24 ;
  LAYER M2 ;
        RECT 5.85 229.18 7.05 229.46 ;
  LAYER M2 ;
        RECT 6.28 234.64 7.48 234.92 ;
  LAYER M2 ;
        RECT 6.28 238.84 7.48 239.12 ;
  LAYER M2 ;
        RECT 5.85 235.06 7.05 235.34 ;
  LAYER M2 ;
        RECT 6.28 240.52 7.48 240.8 ;
  LAYER M2 ;
        RECT 6.28 244.72 7.48 245 ;
  LAYER M2 ;
        RECT 5.85 240.94 7.05 241.22 ;
  LAYER M2 ;
        RECT 6.28 246.4 7.48 246.68 ;
  LAYER M2 ;
        RECT 6.28 250.6 7.48 250.88 ;
  LAYER M2 ;
        RECT 5.85 246.82 7.05 247.1 ;
  LAYER M2 ;
        RECT 6.28 252.28 7.48 252.56 ;
  LAYER M2 ;
        RECT 6.28 256.48 7.48 256.76 ;
  LAYER M2 ;
        RECT 5.85 252.7 7.05 252.98 ;
  LAYER M2 ;
        RECT 6.28 258.16 7.48 258.44 ;
  LAYER M2 ;
        RECT 6.28 262.36 7.48 262.64 ;
  LAYER M2 ;
        RECT 5.85 258.58 7.05 258.86 ;
  LAYER M2 ;
        RECT 6.28 264.04 7.48 264.32 ;
  LAYER M2 ;
        RECT 6.28 268.24 7.48 268.52 ;
  LAYER M2 ;
        RECT 5.85 264.46 7.05 264.74 ;
  LAYER M2 ;
        RECT 6.28 269.92 7.48 270.2 ;
  LAYER M2 ;
        RECT 6.28 274.12 7.48 274.4 ;
  LAYER M2 ;
        RECT 5.85 270.34 7.05 270.62 ;
  LAYER M2 ;
        RECT 6.28 275.8 7.48 276.08 ;
  LAYER M2 ;
        RECT 6.28 280 7.48 280.28 ;
  LAYER M2 ;
        RECT 5.85 276.22 7.05 276.5 ;
  LAYER M2 ;
        RECT 6.28 281.68 7.48 281.96 ;
  LAYER M2 ;
        RECT 6.28 285.88 7.48 286.16 ;
  LAYER M2 ;
        RECT 5.85 282.1 7.05 282.38 ;
  LAYER M2 ;
        RECT 6.28 287.56 7.48 287.84 ;
  LAYER M2 ;
        RECT 6.28 291.76 7.48 292.04 ;
  LAYER M2 ;
        RECT 5.85 287.98 7.05 288.26 ;
  LAYER M2 ;
        RECT 6.28 293.44 7.48 293.72 ;
  LAYER M2 ;
        RECT 6.28 297.64 7.48 297.92 ;
  LAYER M2 ;
        RECT 5.85 293.86 7.05 294.14 ;
  LAYER M2 ;
        RECT 6.28 299.32 7.48 299.6 ;
  LAYER M2 ;
        RECT 6.28 303.52 7.48 303.8 ;
  LAYER M2 ;
        RECT 5.85 299.74 7.05 300.02 ;
  LAYER M2 ;
        RECT 6.28 305.2 7.48 305.48 ;
  LAYER M2 ;
        RECT 6.28 309.4 7.48 309.68 ;
  LAYER M2 ;
        RECT 5.85 305.62 7.05 305.9 ;
  LAYER M2 ;
        RECT 6.28 311.08 7.48 311.36 ;
  LAYER M2 ;
        RECT 6.28 315.28 7.48 315.56 ;
  LAYER M2 ;
        RECT 5.85 311.5 7.05 311.78 ;
  LAYER M2 ;
        RECT 6.28 316.96 7.48 317.24 ;
  LAYER M2 ;
        RECT 6.28 321.16 7.48 321.44 ;
  LAYER M2 ;
        RECT 5.85 317.38 7.05 317.66 ;
  LAYER M2 ;
        RECT 6.28 322.84 7.48 323.12 ;
  LAYER M2 ;
        RECT 6.28 327.04 7.48 327.32 ;
  LAYER M2 ;
        RECT 5.85 323.26 7.05 323.54 ;
  LAYER M2 ;
        RECT 6.28 328.72 7.48 329 ;
  LAYER M2 ;
        RECT 6.28 332.92 7.48 333.2 ;
  LAYER M2 ;
        RECT 5.85 329.14 7.05 329.42 ;
  LAYER M2 ;
        RECT 6.28 334.6 7.48 334.88 ;
  LAYER M2 ;
        RECT 6.28 338.8 7.48 339.08 ;
  LAYER M2 ;
        RECT 5.85 335.02 7.05 335.3 ;
  LAYER M2 ;
        RECT 6.28 340.48 7.48 340.76 ;
  LAYER M2 ;
        RECT 6.28 344.68 7.48 344.96 ;
  LAYER M2 ;
        RECT 5.85 340.9 7.05 341.18 ;
  LAYER M2 ;
        RECT 6.28 346.36 7.48 346.64 ;
  LAYER M2 ;
        RECT 6.28 350.56 7.48 350.84 ;
  LAYER M2 ;
        RECT 5.85 346.78 7.05 347.06 ;
  LAYER M2 ;
        RECT 6.28 352.24 7.48 352.52 ;
  LAYER M2 ;
        RECT 6.28 356.44 7.48 356.72 ;
  LAYER M2 ;
        RECT 5.85 352.66 7.05 352.94 ;
  LAYER M2 ;
        RECT 6.28 358.12 7.48 358.4 ;
  LAYER M2 ;
        RECT 6.28 362.32 7.48 362.6 ;
  LAYER M2 ;
        RECT 5.85 358.54 7.05 358.82 ;
  LAYER M2 ;
        RECT 6.28 364 7.48 364.28 ;
  LAYER M2 ;
        RECT 6.28 368.2 7.48 368.48 ;
  LAYER M2 ;
        RECT 5.85 364.42 7.05 364.7 ;
  LAYER M2 ;
        RECT 6.28 369.88 7.48 370.16 ;
  LAYER M2 ;
        RECT 6.28 374.08 7.48 374.36 ;
  LAYER M2 ;
        RECT 5.85 370.3 7.05 370.58 ;
  LAYER M2 ;
        RECT 6.28 375.76 7.48 376.04 ;
  LAYER M2 ;
        RECT 6.28 379.96 7.48 380.24 ;
  LAYER M2 ;
        RECT 5.85 376.18 7.05 376.46 ;
  LAYER M2 ;
        RECT 6.28 381.64 7.48 381.92 ;
  LAYER M2 ;
        RECT 6.28 385.84 7.48 386.12 ;
  LAYER M2 ;
        RECT 5.85 382.06 7.05 382.34 ;
  LAYER M2 ;
        RECT 6.28 387.52 7.48 387.8 ;
  LAYER M2 ;
        RECT 6.28 391.72 7.48 392 ;
  LAYER M2 ;
        RECT 5.85 387.94 7.05 388.22 ;
  LAYER M2 ;
        RECT 6.28 393.4 7.48 393.68 ;
  LAYER M2 ;
        RECT 6.28 397.6 7.48 397.88 ;
  LAYER M2 ;
        RECT 5.85 393.82 7.05 394.1 ;
  LAYER M2 ;
        RECT 6.28 399.28 7.48 399.56 ;
  LAYER M2 ;
        RECT 6.28 403.48 7.48 403.76 ;
  LAYER M2 ;
        RECT 5.85 399.7 7.05 399.98 ;
  LAYER M2 ;
        RECT 6.28 405.16 7.48 405.44 ;
  LAYER M2 ;
        RECT 6.28 409.36 7.48 409.64 ;
  LAYER M2 ;
        RECT 5.85 405.58 7.05 405.86 ;
  LAYER M2 ;
        RECT 6.28 411.04 7.48 411.32 ;
  LAYER M2 ;
        RECT 6.28 415.24 7.48 415.52 ;
  LAYER M2 ;
        RECT 5.85 411.46 7.05 411.74 ;
  LAYER M2 ;
        RECT 6.28 416.92 7.48 417.2 ;
  LAYER M2 ;
        RECT 6.28 421.12 7.48 421.4 ;
  LAYER M2 ;
        RECT 5.85 417.34 7.05 417.62 ;
  LAYER M2 ;
        RECT 6.28 422.8 7.48 423.08 ;
  LAYER M2 ;
        RECT 6.28 427 7.48 427.28 ;
  LAYER M2 ;
        RECT 5.85 423.22 7.05 423.5 ;
  LAYER M2 ;
        RECT 6.28 428.68 7.48 428.96 ;
  LAYER M2 ;
        RECT 6.28 432.88 7.48 433.16 ;
  LAYER M2 ;
        RECT 5.85 429.1 7.05 429.38 ;
  LAYER M2 ;
        RECT 6.28 434.56 7.48 434.84 ;
  LAYER M2 ;
        RECT 6.28 438.76 7.48 439.04 ;
  LAYER M2 ;
        RECT 5.85 434.98 7.05 435.26 ;
  LAYER M2 ;
        RECT 6.28 440.44 7.48 440.72 ;
  LAYER M2 ;
        RECT 6.28 444.64 7.48 444.92 ;
  LAYER M2 ;
        RECT 5.85 440.86 7.05 441.14 ;
  LAYER M2 ;
        RECT 6.28 446.32 7.48 446.6 ;
  LAYER M2 ;
        RECT 6.28 450.52 7.48 450.8 ;
  LAYER M2 ;
        RECT 5.85 446.74 7.05 447.02 ;
  LAYER M2 ;
        RECT 6.28 452.2 7.48 452.48 ;
  LAYER M2 ;
        RECT 6.28 456.4 7.48 456.68 ;
  LAYER M2 ;
        RECT 5.85 452.62 7.05 452.9 ;
  LAYER M2 ;
        RECT 6.28 458.08 7.48 458.36 ;
  LAYER M2 ;
        RECT 6.28 462.28 7.48 462.56 ;
  LAYER M2 ;
        RECT 5.85 458.5 7.05 458.78 ;
  LAYER M2 ;
        RECT 6.28 463.96 7.48 464.24 ;
  LAYER M2 ;
        RECT 6.28 468.16 7.48 468.44 ;
  LAYER M2 ;
        RECT 5.85 464.38 7.05 464.66 ;
  LAYER M2 ;
        RECT 6.28 469.84 7.48 470.12 ;
  LAYER M2 ;
        RECT 6.28 474.04 7.48 474.32 ;
  LAYER M2 ;
        RECT 5.85 470.26 7.05 470.54 ;
  LAYER M2 ;
        RECT 6.28 475.72 7.48 476 ;
  LAYER M2 ;
        RECT 6.28 479.92 7.48 480.2 ;
  LAYER M2 ;
        RECT 5.85 476.14 7.05 476.42 ;
  LAYER M2 ;
        RECT 5.85 482.02 7.05 482.3 ;
  LAYER M3 ;
        RECT 6.74 64.1 7.02 476.02 ;
  LAYER M3 ;
        RECT 6.31 68.3 6.59 480.22 ;
  LAYER M3 ;
        RECT 5.88 64.52 6.16 482.32 ;
  LAYER M1 ;
        RECT 3.745 33.095 3.995 36.625 ;
  LAYER M1 ;
        RECT 3.745 31.835 3.995 32.845 ;
  LAYER M1 ;
        RECT 3.745 27.215 3.995 30.745 ;
  LAYER M1 ;
        RECT 3.745 25.955 3.995 26.965 ;
  LAYER M1 ;
        RECT 3.745 21.335 3.995 24.865 ;
  LAYER M1 ;
        RECT 3.745 20.075 3.995 21.085 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 18.985 ;
  LAYER M1 ;
        RECT 3.745 14.195 3.995 15.205 ;
  LAYER M1 ;
        RECT 3.745 9.575 3.995 13.105 ;
  LAYER M1 ;
        RECT 3.745 8.315 3.995 9.325 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 33.095 4.425 36.625 ;
  LAYER M1 ;
        RECT 4.175 27.215 4.425 30.745 ;
  LAYER M1 ;
        RECT 4.175 21.335 4.425 24.865 ;
  LAYER M1 ;
        RECT 4.175 15.455 4.425 18.985 ;
  LAYER M1 ;
        RECT 4.175 9.575 4.425 13.105 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 33.095 3.565 36.625 ;
  LAYER M1 ;
        RECT 3.315 27.215 3.565 30.745 ;
  LAYER M1 ;
        RECT 3.315 21.335 3.565 24.865 ;
  LAYER M1 ;
        RECT 3.315 15.455 3.565 18.985 ;
  LAYER M1 ;
        RECT 3.315 9.575 3.565 13.105 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 2.885 33.095 3.135 36.625 ;
  LAYER M1 ;
        RECT 2.885 31.835 3.135 32.845 ;
  LAYER M1 ;
        RECT 2.885 27.215 3.135 30.745 ;
  LAYER M1 ;
        RECT 2.885 25.955 3.135 26.965 ;
  LAYER M1 ;
        RECT 2.885 21.335 3.135 24.865 ;
  LAYER M1 ;
        RECT 2.885 20.075 3.135 21.085 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 18.985 ;
  LAYER M1 ;
        RECT 2.885 14.195 3.135 15.205 ;
  LAYER M1 ;
        RECT 2.885 9.575 3.135 13.105 ;
  LAYER M1 ;
        RECT 2.885 8.315 3.135 9.325 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 2.455 33.095 2.705 36.625 ;
  LAYER M1 ;
        RECT 2.455 27.215 2.705 30.745 ;
  LAYER M1 ;
        RECT 2.455 21.335 2.705 24.865 ;
  LAYER M1 ;
        RECT 2.455 15.455 2.705 18.985 ;
  LAYER M1 ;
        RECT 2.455 9.575 2.705 13.105 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.025 33.095 2.275 36.625 ;
  LAYER M1 ;
        RECT 2.025 31.835 2.275 32.845 ;
  LAYER M1 ;
        RECT 2.025 27.215 2.275 30.745 ;
  LAYER M1 ;
        RECT 2.025 25.955 2.275 26.965 ;
  LAYER M1 ;
        RECT 2.025 21.335 2.275 24.865 ;
  LAYER M1 ;
        RECT 2.025 20.075 2.275 21.085 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 18.985 ;
  LAYER M1 ;
        RECT 2.025 14.195 2.275 15.205 ;
  LAYER M1 ;
        RECT 2.025 9.575 2.275 13.105 ;
  LAYER M1 ;
        RECT 2.025 8.315 2.275 9.325 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 1.595 33.095 1.845 36.625 ;
  LAYER M1 ;
        RECT 1.595 27.215 1.845 30.745 ;
  LAYER M1 ;
        RECT 1.595 21.335 1.845 24.865 ;
  LAYER M1 ;
        RECT 1.595 15.455 1.845 18.985 ;
  LAYER M1 ;
        RECT 1.595 9.575 1.845 13.105 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 1.98 36.4 4.04 36.68 ;
  LAYER M2 ;
        RECT 1.98 32.2 4.04 32.48 ;
  LAYER M2 ;
        RECT 1.55 35.98 4.47 36.26 ;
  LAYER M2 ;
        RECT 1.98 30.52 4.04 30.8 ;
  LAYER M2 ;
        RECT 1.98 26.32 4.04 26.6 ;
  LAYER M2 ;
        RECT 1.55 30.1 4.47 30.38 ;
  LAYER M2 ;
        RECT 1.98 24.64 4.04 24.92 ;
  LAYER M2 ;
        RECT 1.98 20.44 4.04 20.72 ;
  LAYER M2 ;
        RECT 1.55 24.22 4.47 24.5 ;
  LAYER M2 ;
        RECT 1.98 18.76 4.04 19.04 ;
  LAYER M2 ;
        RECT 1.98 14.56 4.04 14.84 ;
  LAYER M2 ;
        RECT 1.55 18.34 4.47 18.62 ;
  LAYER M2 ;
        RECT 1.98 12.88 4.04 13.16 ;
  LAYER M2 ;
        RECT 1.98 8.68 4.04 8.96 ;
  LAYER M2 ;
        RECT 1.55 12.46 4.47 12.74 ;
  LAYER M2 ;
        RECT 1.98 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 1.98 2.8 4.04 3.08 ;
  LAYER M2 ;
        RECT 1.55 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 1.98 0.7 4.04 0.98 ;
  LAYER M3 ;
        RECT 3.3 6.98 3.58 36.7 ;
  LAYER M3 ;
        RECT 2.87 2.78 3.15 32.5 ;
  LAYER M3 ;
        RECT 2.44 0.68 2.72 36.28 ;
  LAYER M1 ;
        RECT 1.165 208.655 1.415 212.185 ;
  LAYER M1 ;
        RECT 1.165 207.395 1.415 208.405 ;
  LAYER M1 ;
        RECT 1.165 202.775 1.415 206.305 ;
  LAYER M1 ;
        RECT 1.165 201.515 1.415 202.525 ;
  LAYER M1 ;
        RECT 1.165 196.895 1.415 200.425 ;
  LAYER M1 ;
        RECT 1.165 195.635 1.415 196.645 ;
  LAYER M1 ;
        RECT 1.165 191.015 1.415 194.545 ;
  LAYER M1 ;
        RECT 1.165 189.755 1.415 190.765 ;
  LAYER M1 ;
        RECT 1.165 185.135 1.415 188.665 ;
  LAYER M1 ;
        RECT 1.165 183.875 1.415 184.885 ;
  LAYER M1 ;
        RECT 1.165 179.255 1.415 182.785 ;
  LAYER M1 ;
        RECT 1.165 177.995 1.415 179.005 ;
  LAYER M1 ;
        RECT 1.165 173.375 1.415 176.905 ;
  LAYER M1 ;
        RECT 1.165 172.115 1.415 173.125 ;
  LAYER M1 ;
        RECT 1.165 167.495 1.415 171.025 ;
  LAYER M1 ;
        RECT 1.165 166.235 1.415 167.245 ;
  LAYER M1 ;
        RECT 1.165 161.615 1.415 165.145 ;
  LAYER M1 ;
        RECT 1.165 160.355 1.415 161.365 ;
  LAYER M1 ;
        RECT 1.165 155.735 1.415 159.265 ;
  LAYER M1 ;
        RECT 1.165 154.475 1.415 155.485 ;
  LAYER M1 ;
        RECT 1.165 149.855 1.415 153.385 ;
  LAYER M1 ;
        RECT 1.165 148.595 1.415 149.605 ;
  LAYER M1 ;
        RECT 1.165 143.975 1.415 147.505 ;
  LAYER M1 ;
        RECT 1.165 142.715 1.415 143.725 ;
  LAYER M1 ;
        RECT 1.165 138.095 1.415 141.625 ;
  LAYER M1 ;
        RECT 1.165 136.835 1.415 137.845 ;
  LAYER M1 ;
        RECT 1.165 132.215 1.415 135.745 ;
  LAYER M1 ;
        RECT 1.165 130.955 1.415 131.965 ;
  LAYER M1 ;
        RECT 1.165 126.335 1.415 129.865 ;
  LAYER M1 ;
        RECT 1.165 125.075 1.415 126.085 ;
  LAYER M1 ;
        RECT 1.165 120.455 1.415 123.985 ;
  LAYER M1 ;
        RECT 1.165 119.195 1.415 120.205 ;
  LAYER M1 ;
        RECT 1.165 114.575 1.415 118.105 ;
  LAYER M1 ;
        RECT 1.165 113.315 1.415 114.325 ;
  LAYER M1 ;
        RECT 1.165 108.695 1.415 112.225 ;
  LAYER M1 ;
        RECT 1.165 107.435 1.415 108.445 ;
  LAYER M1 ;
        RECT 1.165 102.815 1.415 106.345 ;
  LAYER M1 ;
        RECT 1.165 101.555 1.415 102.565 ;
  LAYER M1 ;
        RECT 1.165 96.935 1.415 100.465 ;
  LAYER M1 ;
        RECT 1.165 95.675 1.415 96.685 ;
  LAYER M1 ;
        RECT 1.165 91.055 1.415 94.585 ;
  LAYER M1 ;
        RECT 1.165 89.795 1.415 90.805 ;
  LAYER M1 ;
        RECT 1.165 85.175 1.415 88.705 ;
  LAYER M1 ;
        RECT 1.165 83.915 1.415 84.925 ;
  LAYER M1 ;
        RECT 1.165 79.295 1.415 82.825 ;
  LAYER M1 ;
        RECT 1.165 78.035 1.415 79.045 ;
  LAYER M1 ;
        RECT 1.165 73.415 1.415 76.945 ;
  LAYER M1 ;
        RECT 1.165 72.155 1.415 73.165 ;
  LAYER M1 ;
        RECT 1.165 67.535 1.415 71.065 ;
  LAYER M1 ;
        RECT 1.165 66.275 1.415 67.285 ;
  LAYER M1 ;
        RECT 1.165 64.175 1.415 65.185 ;
  LAYER M1 ;
        RECT 1.595 208.655 1.845 212.185 ;
  LAYER M1 ;
        RECT 1.595 202.775 1.845 206.305 ;
  LAYER M1 ;
        RECT 1.595 196.895 1.845 200.425 ;
  LAYER M1 ;
        RECT 1.595 191.015 1.845 194.545 ;
  LAYER M1 ;
        RECT 1.595 185.135 1.845 188.665 ;
  LAYER M1 ;
        RECT 1.595 179.255 1.845 182.785 ;
  LAYER M1 ;
        RECT 1.595 173.375 1.845 176.905 ;
  LAYER M1 ;
        RECT 1.595 167.495 1.845 171.025 ;
  LAYER M1 ;
        RECT 1.595 161.615 1.845 165.145 ;
  LAYER M1 ;
        RECT 1.595 155.735 1.845 159.265 ;
  LAYER M1 ;
        RECT 1.595 149.855 1.845 153.385 ;
  LAYER M1 ;
        RECT 1.595 143.975 1.845 147.505 ;
  LAYER M1 ;
        RECT 1.595 138.095 1.845 141.625 ;
  LAYER M1 ;
        RECT 1.595 132.215 1.845 135.745 ;
  LAYER M1 ;
        RECT 1.595 126.335 1.845 129.865 ;
  LAYER M1 ;
        RECT 1.595 120.455 1.845 123.985 ;
  LAYER M1 ;
        RECT 1.595 114.575 1.845 118.105 ;
  LAYER M1 ;
        RECT 1.595 108.695 1.845 112.225 ;
  LAYER M1 ;
        RECT 1.595 102.815 1.845 106.345 ;
  LAYER M1 ;
        RECT 1.595 96.935 1.845 100.465 ;
  LAYER M1 ;
        RECT 1.595 91.055 1.845 94.585 ;
  LAYER M1 ;
        RECT 1.595 85.175 1.845 88.705 ;
  LAYER M1 ;
        RECT 1.595 79.295 1.845 82.825 ;
  LAYER M1 ;
        RECT 1.595 73.415 1.845 76.945 ;
  LAYER M1 ;
        RECT 1.595 67.535 1.845 71.065 ;
  LAYER M1 ;
        RECT 0.735 208.655 0.985 212.185 ;
  LAYER M1 ;
        RECT 0.735 202.775 0.985 206.305 ;
  LAYER M1 ;
        RECT 0.735 196.895 0.985 200.425 ;
  LAYER M1 ;
        RECT 0.735 191.015 0.985 194.545 ;
  LAYER M1 ;
        RECT 0.735 185.135 0.985 188.665 ;
  LAYER M1 ;
        RECT 0.735 179.255 0.985 182.785 ;
  LAYER M1 ;
        RECT 0.735 173.375 0.985 176.905 ;
  LAYER M1 ;
        RECT 0.735 167.495 0.985 171.025 ;
  LAYER M1 ;
        RECT 0.735 161.615 0.985 165.145 ;
  LAYER M1 ;
        RECT 0.735 155.735 0.985 159.265 ;
  LAYER M1 ;
        RECT 0.735 149.855 0.985 153.385 ;
  LAYER M1 ;
        RECT 0.735 143.975 0.985 147.505 ;
  LAYER M1 ;
        RECT 0.735 138.095 0.985 141.625 ;
  LAYER M1 ;
        RECT 0.735 132.215 0.985 135.745 ;
  LAYER M1 ;
        RECT 0.735 126.335 0.985 129.865 ;
  LAYER M1 ;
        RECT 0.735 120.455 0.985 123.985 ;
  LAYER M1 ;
        RECT 0.735 114.575 0.985 118.105 ;
  LAYER M1 ;
        RECT 0.735 108.695 0.985 112.225 ;
  LAYER M1 ;
        RECT 0.735 102.815 0.985 106.345 ;
  LAYER M1 ;
        RECT 0.735 96.935 0.985 100.465 ;
  LAYER M1 ;
        RECT 0.735 91.055 0.985 94.585 ;
  LAYER M1 ;
        RECT 0.735 85.175 0.985 88.705 ;
  LAYER M1 ;
        RECT 0.735 79.295 0.985 82.825 ;
  LAYER M1 ;
        RECT 0.735 73.415 0.985 76.945 ;
  LAYER M1 ;
        RECT 0.735 67.535 0.985 71.065 ;
  LAYER M2 ;
        RECT 1.12 211.96 2.32 212.24 ;
  LAYER M2 ;
        RECT 1.12 207.76 2.32 208.04 ;
  LAYER M2 ;
        RECT 0.69 211.54 1.89 211.82 ;
  LAYER M2 ;
        RECT 1.12 206.08 2.32 206.36 ;
  LAYER M2 ;
        RECT 1.12 201.88 2.32 202.16 ;
  LAYER M2 ;
        RECT 0.69 205.66 1.89 205.94 ;
  LAYER M2 ;
        RECT 1.12 200.2 2.32 200.48 ;
  LAYER M2 ;
        RECT 1.12 196 2.32 196.28 ;
  LAYER M2 ;
        RECT 0.69 199.78 1.89 200.06 ;
  LAYER M2 ;
        RECT 1.12 194.32 2.32 194.6 ;
  LAYER M2 ;
        RECT 1.12 190.12 2.32 190.4 ;
  LAYER M2 ;
        RECT 0.69 193.9 1.89 194.18 ;
  LAYER M2 ;
        RECT 1.12 188.44 2.32 188.72 ;
  LAYER M2 ;
        RECT 1.12 184.24 2.32 184.52 ;
  LAYER M2 ;
        RECT 0.69 188.02 1.89 188.3 ;
  LAYER M2 ;
        RECT 1.12 182.56 2.32 182.84 ;
  LAYER M2 ;
        RECT 1.12 178.36 2.32 178.64 ;
  LAYER M2 ;
        RECT 0.69 182.14 1.89 182.42 ;
  LAYER M2 ;
        RECT 1.12 176.68 2.32 176.96 ;
  LAYER M2 ;
        RECT 1.12 172.48 2.32 172.76 ;
  LAYER M2 ;
        RECT 0.69 176.26 1.89 176.54 ;
  LAYER M2 ;
        RECT 1.12 170.8 2.32 171.08 ;
  LAYER M2 ;
        RECT 1.12 166.6 2.32 166.88 ;
  LAYER M2 ;
        RECT 0.69 170.38 1.89 170.66 ;
  LAYER M2 ;
        RECT 1.12 164.92 2.32 165.2 ;
  LAYER M2 ;
        RECT 1.12 160.72 2.32 161 ;
  LAYER M2 ;
        RECT 0.69 164.5 1.89 164.78 ;
  LAYER M2 ;
        RECT 1.12 159.04 2.32 159.32 ;
  LAYER M2 ;
        RECT 1.12 154.84 2.32 155.12 ;
  LAYER M2 ;
        RECT 0.69 158.62 1.89 158.9 ;
  LAYER M2 ;
        RECT 1.12 153.16 2.32 153.44 ;
  LAYER M2 ;
        RECT 1.12 148.96 2.32 149.24 ;
  LAYER M2 ;
        RECT 0.69 152.74 1.89 153.02 ;
  LAYER M2 ;
        RECT 1.12 147.28 2.32 147.56 ;
  LAYER M2 ;
        RECT 1.12 143.08 2.32 143.36 ;
  LAYER M2 ;
        RECT 0.69 146.86 1.89 147.14 ;
  LAYER M2 ;
        RECT 1.12 141.4 2.32 141.68 ;
  LAYER M2 ;
        RECT 1.12 137.2 2.32 137.48 ;
  LAYER M2 ;
        RECT 0.69 140.98 1.89 141.26 ;
  LAYER M2 ;
        RECT 1.12 135.52 2.32 135.8 ;
  LAYER M2 ;
        RECT 1.12 131.32 2.32 131.6 ;
  LAYER M2 ;
        RECT 0.69 135.1 1.89 135.38 ;
  LAYER M2 ;
        RECT 1.12 129.64 2.32 129.92 ;
  LAYER M2 ;
        RECT 1.12 125.44 2.32 125.72 ;
  LAYER M2 ;
        RECT 0.69 129.22 1.89 129.5 ;
  LAYER M2 ;
        RECT 1.12 123.76 2.32 124.04 ;
  LAYER M2 ;
        RECT 1.12 119.56 2.32 119.84 ;
  LAYER M2 ;
        RECT 0.69 123.34 1.89 123.62 ;
  LAYER M2 ;
        RECT 1.12 117.88 2.32 118.16 ;
  LAYER M2 ;
        RECT 1.12 113.68 2.32 113.96 ;
  LAYER M2 ;
        RECT 0.69 117.46 1.89 117.74 ;
  LAYER M2 ;
        RECT 1.12 112 2.32 112.28 ;
  LAYER M2 ;
        RECT 1.12 107.8 2.32 108.08 ;
  LAYER M2 ;
        RECT 0.69 111.58 1.89 111.86 ;
  LAYER M2 ;
        RECT 1.12 106.12 2.32 106.4 ;
  LAYER M2 ;
        RECT 1.12 101.92 2.32 102.2 ;
  LAYER M2 ;
        RECT 0.69 105.7 1.89 105.98 ;
  LAYER M2 ;
        RECT 1.12 100.24 2.32 100.52 ;
  LAYER M2 ;
        RECT 1.12 96.04 2.32 96.32 ;
  LAYER M2 ;
        RECT 0.69 99.82 1.89 100.1 ;
  LAYER M2 ;
        RECT 1.12 94.36 2.32 94.64 ;
  LAYER M2 ;
        RECT 1.12 90.16 2.32 90.44 ;
  LAYER M2 ;
        RECT 0.69 93.94 1.89 94.22 ;
  LAYER M2 ;
        RECT 1.12 88.48 2.32 88.76 ;
  LAYER M2 ;
        RECT 1.12 84.28 2.32 84.56 ;
  LAYER M2 ;
        RECT 0.69 88.06 1.89 88.34 ;
  LAYER M2 ;
        RECT 1.12 82.6 2.32 82.88 ;
  LAYER M2 ;
        RECT 1.12 78.4 2.32 78.68 ;
  LAYER M2 ;
        RECT 0.69 82.18 1.89 82.46 ;
  LAYER M2 ;
        RECT 1.12 76.72 2.32 77 ;
  LAYER M2 ;
        RECT 1.12 72.52 2.32 72.8 ;
  LAYER M2 ;
        RECT 0.69 76.3 1.89 76.58 ;
  LAYER M2 ;
        RECT 1.12 70.84 2.32 71.12 ;
  LAYER M2 ;
        RECT 1.12 66.64 2.32 66.92 ;
  LAYER M2 ;
        RECT 0.69 70.42 1.89 70.7 ;
  LAYER M2 ;
        RECT 0.69 64.54 1.89 64.82 ;
  LAYER M3 ;
        RECT 1.58 70.82 1.86 212.26 ;
  LAYER M3 ;
        RECT 1.15 66.62 1.43 208.06 ;
  LAYER M3 ;
        RECT 0.72 64.52 1 211.84 ;
  LAYER M1 ;
        RECT 8.905 208.655 9.155 212.185 ;
  LAYER M1 ;
        RECT 8.905 207.395 9.155 208.405 ;
  LAYER M1 ;
        RECT 8.905 202.775 9.155 206.305 ;
  LAYER M1 ;
        RECT 8.905 201.515 9.155 202.525 ;
  LAYER M1 ;
        RECT 8.905 196.895 9.155 200.425 ;
  LAYER M1 ;
        RECT 8.905 195.635 9.155 196.645 ;
  LAYER M1 ;
        RECT 8.905 191.015 9.155 194.545 ;
  LAYER M1 ;
        RECT 8.905 189.755 9.155 190.765 ;
  LAYER M1 ;
        RECT 8.905 185.135 9.155 188.665 ;
  LAYER M1 ;
        RECT 8.905 183.875 9.155 184.885 ;
  LAYER M1 ;
        RECT 8.905 179.255 9.155 182.785 ;
  LAYER M1 ;
        RECT 8.905 177.995 9.155 179.005 ;
  LAYER M1 ;
        RECT 8.905 173.375 9.155 176.905 ;
  LAYER M1 ;
        RECT 8.905 172.115 9.155 173.125 ;
  LAYER M1 ;
        RECT 8.905 167.495 9.155 171.025 ;
  LAYER M1 ;
        RECT 8.905 166.235 9.155 167.245 ;
  LAYER M1 ;
        RECT 8.905 161.615 9.155 165.145 ;
  LAYER M1 ;
        RECT 8.905 160.355 9.155 161.365 ;
  LAYER M1 ;
        RECT 8.905 155.735 9.155 159.265 ;
  LAYER M1 ;
        RECT 8.905 154.475 9.155 155.485 ;
  LAYER M1 ;
        RECT 8.905 149.855 9.155 153.385 ;
  LAYER M1 ;
        RECT 8.905 148.595 9.155 149.605 ;
  LAYER M1 ;
        RECT 8.905 143.975 9.155 147.505 ;
  LAYER M1 ;
        RECT 8.905 142.715 9.155 143.725 ;
  LAYER M1 ;
        RECT 8.905 138.095 9.155 141.625 ;
  LAYER M1 ;
        RECT 8.905 136.835 9.155 137.845 ;
  LAYER M1 ;
        RECT 8.905 132.215 9.155 135.745 ;
  LAYER M1 ;
        RECT 8.905 130.955 9.155 131.965 ;
  LAYER M1 ;
        RECT 8.905 126.335 9.155 129.865 ;
  LAYER M1 ;
        RECT 8.905 125.075 9.155 126.085 ;
  LAYER M1 ;
        RECT 8.905 120.455 9.155 123.985 ;
  LAYER M1 ;
        RECT 8.905 119.195 9.155 120.205 ;
  LAYER M1 ;
        RECT 8.905 114.575 9.155 118.105 ;
  LAYER M1 ;
        RECT 8.905 113.315 9.155 114.325 ;
  LAYER M1 ;
        RECT 8.905 108.695 9.155 112.225 ;
  LAYER M1 ;
        RECT 8.905 107.435 9.155 108.445 ;
  LAYER M1 ;
        RECT 8.905 102.815 9.155 106.345 ;
  LAYER M1 ;
        RECT 8.905 101.555 9.155 102.565 ;
  LAYER M1 ;
        RECT 8.905 96.935 9.155 100.465 ;
  LAYER M1 ;
        RECT 8.905 95.675 9.155 96.685 ;
  LAYER M1 ;
        RECT 8.905 91.055 9.155 94.585 ;
  LAYER M1 ;
        RECT 8.905 89.795 9.155 90.805 ;
  LAYER M1 ;
        RECT 8.905 85.175 9.155 88.705 ;
  LAYER M1 ;
        RECT 8.905 83.915 9.155 84.925 ;
  LAYER M1 ;
        RECT 8.905 79.295 9.155 82.825 ;
  LAYER M1 ;
        RECT 8.905 78.035 9.155 79.045 ;
  LAYER M1 ;
        RECT 8.905 73.415 9.155 76.945 ;
  LAYER M1 ;
        RECT 8.905 72.155 9.155 73.165 ;
  LAYER M1 ;
        RECT 8.905 67.535 9.155 71.065 ;
  LAYER M1 ;
        RECT 8.905 66.275 9.155 67.285 ;
  LAYER M1 ;
        RECT 8.905 64.175 9.155 65.185 ;
  LAYER M1 ;
        RECT 8.475 208.655 8.725 212.185 ;
  LAYER M1 ;
        RECT 8.475 202.775 8.725 206.305 ;
  LAYER M1 ;
        RECT 8.475 196.895 8.725 200.425 ;
  LAYER M1 ;
        RECT 8.475 191.015 8.725 194.545 ;
  LAYER M1 ;
        RECT 8.475 185.135 8.725 188.665 ;
  LAYER M1 ;
        RECT 8.475 179.255 8.725 182.785 ;
  LAYER M1 ;
        RECT 8.475 173.375 8.725 176.905 ;
  LAYER M1 ;
        RECT 8.475 167.495 8.725 171.025 ;
  LAYER M1 ;
        RECT 8.475 161.615 8.725 165.145 ;
  LAYER M1 ;
        RECT 8.475 155.735 8.725 159.265 ;
  LAYER M1 ;
        RECT 8.475 149.855 8.725 153.385 ;
  LAYER M1 ;
        RECT 8.475 143.975 8.725 147.505 ;
  LAYER M1 ;
        RECT 8.475 138.095 8.725 141.625 ;
  LAYER M1 ;
        RECT 8.475 132.215 8.725 135.745 ;
  LAYER M1 ;
        RECT 8.475 126.335 8.725 129.865 ;
  LAYER M1 ;
        RECT 8.475 120.455 8.725 123.985 ;
  LAYER M1 ;
        RECT 8.475 114.575 8.725 118.105 ;
  LAYER M1 ;
        RECT 8.475 108.695 8.725 112.225 ;
  LAYER M1 ;
        RECT 8.475 102.815 8.725 106.345 ;
  LAYER M1 ;
        RECT 8.475 96.935 8.725 100.465 ;
  LAYER M1 ;
        RECT 8.475 91.055 8.725 94.585 ;
  LAYER M1 ;
        RECT 8.475 85.175 8.725 88.705 ;
  LAYER M1 ;
        RECT 8.475 79.295 8.725 82.825 ;
  LAYER M1 ;
        RECT 8.475 73.415 8.725 76.945 ;
  LAYER M1 ;
        RECT 8.475 67.535 8.725 71.065 ;
  LAYER M1 ;
        RECT 9.335 208.655 9.585 212.185 ;
  LAYER M1 ;
        RECT 9.335 202.775 9.585 206.305 ;
  LAYER M1 ;
        RECT 9.335 196.895 9.585 200.425 ;
  LAYER M1 ;
        RECT 9.335 191.015 9.585 194.545 ;
  LAYER M1 ;
        RECT 9.335 185.135 9.585 188.665 ;
  LAYER M1 ;
        RECT 9.335 179.255 9.585 182.785 ;
  LAYER M1 ;
        RECT 9.335 173.375 9.585 176.905 ;
  LAYER M1 ;
        RECT 9.335 167.495 9.585 171.025 ;
  LAYER M1 ;
        RECT 9.335 161.615 9.585 165.145 ;
  LAYER M1 ;
        RECT 9.335 155.735 9.585 159.265 ;
  LAYER M1 ;
        RECT 9.335 149.855 9.585 153.385 ;
  LAYER M1 ;
        RECT 9.335 143.975 9.585 147.505 ;
  LAYER M1 ;
        RECT 9.335 138.095 9.585 141.625 ;
  LAYER M1 ;
        RECT 9.335 132.215 9.585 135.745 ;
  LAYER M1 ;
        RECT 9.335 126.335 9.585 129.865 ;
  LAYER M1 ;
        RECT 9.335 120.455 9.585 123.985 ;
  LAYER M1 ;
        RECT 9.335 114.575 9.585 118.105 ;
  LAYER M1 ;
        RECT 9.335 108.695 9.585 112.225 ;
  LAYER M1 ;
        RECT 9.335 102.815 9.585 106.345 ;
  LAYER M1 ;
        RECT 9.335 96.935 9.585 100.465 ;
  LAYER M1 ;
        RECT 9.335 91.055 9.585 94.585 ;
  LAYER M1 ;
        RECT 9.335 85.175 9.585 88.705 ;
  LAYER M1 ;
        RECT 9.335 79.295 9.585 82.825 ;
  LAYER M1 ;
        RECT 9.335 73.415 9.585 76.945 ;
  LAYER M1 ;
        RECT 9.335 67.535 9.585 71.065 ;
  LAYER M2 ;
        RECT 8 211.96 9.2 212.24 ;
  LAYER M2 ;
        RECT 8 207.76 9.2 208.04 ;
  LAYER M2 ;
        RECT 8.43 211.54 9.63 211.82 ;
  LAYER M2 ;
        RECT 8 206.08 9.2 206.36 ;
  LAYER M2 ;
        RECT 8 201.88 9.2 202.16 ;
  LAYER M2 ;
        RECT 8.43 205.66 9.63 205.94 ;
  LAYER M2 ;
        RECT 8 200.2 9.2 200.48 ;
  LAYER M2 ;
        RECT 8 196 9.2 196.28 ;
  LAYER M2 ;
        RECT 8.43 199.78 9.63 200.06 ;
  LAYER M2 ;
        RECT 8 194.32 9.2 194.6 ;
  LAYER M2 ;
        RECT 8 190.12 9.2 190.4 ;
  LAYER M2 ;
        RECT 8.43 193.9 9.63 194.18 ;
  LAYER M2 ;
        RECT 8 188.44 9.2 188.72 ;
  LAYER M2 ;
        RECT 8 184.24 9.2 184.52 ;
  LAYER M2 ;
        RECT 8.43 188.02 9.63 188.3 ;
  LAYER M2 ;
        RECT 8 182.56 9.2 182.84 ;
  LAYER M2 ;
        RECT 8 178.36 9.2 178.64 ;
  LAYER M2 ;
        RECT 8.43 182.14 9.63 182.42 ;
  LAYER M2 ;
        RECT 8 176.68 9.2 176.96 ;
  LAYER M2 ;
        RECT 8 172.48 9.2 172.76 ;
  LAYER M2 ;
        RECT 8.43 176.26 9.63 176.54 ;
  LAYER M2 ;
        RECT 8 170.8 9.2 171.08 ;
  LAYER M2 ;
        RECT 8 166.6 9.2 166.88 ;
  LAYER M2 ;
        RECT 8.43 170.38 9.63 170.66 ;
  LAYER M2 ;
        RECT 8 164.92 9.2 165.2 ;
  LAYER M2 ;
        RECT 8 160.72 9.2 161 ;
  LAYER M2 ;
        RECT 8.43 164.5 9.63 164.78 ;
  LAYER M2 ;
        RECT 8 159.04 9.2 159.32 ;
  LAYER M2 ;
        RECT 8 154.84 9.2 155.12 ;
  LAYER M2 ;
        RECT 8.43 158.62 9.63 158.9 ;
  LAYER M2 ;
        RECT 8 153.16 9.2 153.44 ;
  LAYER M2 ;
        RECT 8 148.96 9.2 149.24 ;
  LAYER M2 ;
        RECT 8.43 152.74 9.63 153.02 ;
  LAYER M2 ;
        RECT 8 147.28 9.2 147.56 ;
  LAYER M2 ;
        RECT 8 143.08 9.2 143.36 ;
  LAYER M2 ;
        RECT 8.43 146.86 9.63 147.14 ;
  LAYER M2 ;
        RECT 8 141.4 9.2 141.68 ;
  LAYER M2 ;
        RECT 8 137.2 9.2 137.48 ;
  LAYER M2 ;
        RECT 8.43 140.98 9.63 141.26 ;
  LAYER M2 ;
        RECT 8 135.52 9.2 135.8 ;
  LAYER M2 ;
        RECT 8 131.32 9.2 131.6 ;
  LAYER M2 ;
        RECT 8.43 135.1 9.63 135.38 ;
  LAYER M2 ;
        RECT 8 129.64 9.2 129.92 ;
  LAYER M2 ;
        RECT 8 125.44 9.2 125.72 ;
  LAYER M2 ;
        RECT 8.43 129.22 9.63 129.5 ;
  LAYER M2 ;
        RECT 8 123.76 9.2 124.04 ;
  LAYER M2 ;
        RECT 8 119.56 9.2 119.84 ;
  LAYER M2 ;
        RECT 8.43 123.34 9.63 123.62 ;
  LAYER M2 ;
        RECT 8 117.88 9.2 118.16 ;
  LAYER M2 ;
        RECT 8 113.68 9.2 113.96 ;
  LAYER M2 ;
        RECT 8.43 117.46 9.63 117.74 ;
  LAYER M2 ;
        RECT 8 112 9.2 112.28 ;
  LAYER M2 ;
        RECT 8 107.8 9.2 108.08 ;
  LAYER M2 ;
        RECT 8.43 111.58 9.63 111.86 ;
  LAYER M2 ;
        RECT 8 106.12 9.2 106.4 ;
  LAYER M2 ;
        RECT 8 101.92 9.2 102.2 ;
  LAYER M2 ;
        RECT 8.43 105.7 9.63 105.98 ;
  LAYER M2 ;
        RECT 8 100.24 9.2 100.52 ;
  LAYER M2 ;
        RECT 8 96.04 9.2 96.32 ;
  LAYER M2 ;
        RECT 8.43 99.82 9.63 100.1 ;
  LAYER M2 ;
        RECT 8 94.36 9.2 94.64 ;
  LAYER M2 ;
        RECT 8 90.16 9.2 90.44 ;
  LAYER M2 ;
        RECT 8.43 93.94 9.63 94.22 ;
  LAYER M2 ;
        RECT 8 88.48 9.2 88.76 ;
  LAYER M2 ;
        RECT 8 84.28 9.2 84.56 ;
  LAYER M2 ;
        RECT 8.43 88.06 9.63 88.34 ;
  LAYER M2 ;
        RECT 8 82.6 9.2 82.88 ;
  LAYER M2 ;
        RECT 8 78.4 9.2 78.68 ;
  LAYER M2 ;
        RECT 8.43 82.18 9.63 82.46 ;
  LAYER M2 ;
        RECT 8 76.72 9.2 77 ;
  LAYER M2 ;
        RECT 8 72.52 9.2 72.8 ;
  LAYER M2 ;
        RECT 8.43 76.3 9.63 76.58 ;
  LAYER M2 ;
        RECT 8 70.84 9.2 71.12 ;
  LAYER M2 ;
        RECT 8 66.64 9.2 66.92 ;
  LAYER M2 ;
        RECT 8.43 70.42 9.63 70.7 ;
  LAYER M2 ;
        RECT 8.43 64.54 9.63 64.82 ;
  LAYER M3 ;
        RECT 8.46 70.82 8.74 212.26 ;
  LAYER M3 ;
        RECT 8.89 66.62 9.17 208.06 ;
  LAYER M3 ;
        RECT 9.32 64.52 9.6 211.84 ;
  LAYER M1 ;
        RECT 1.595 52.415 1.845 55.945 ;
  LAYER M1 ;
        RECT 1.595 51.155 1.845 52.165 ;
  LAYER M1 ;
        RECT 1.595 46.535 1.845 50.065 ;
  LAYER M1 ;
        RECT 1.595 45.275 1.845 46.285 ;
  LAYER M1 ;
        RECT 1.595 40.655 1.845 44.185 ;
  LAYER M1 ;
        RECT 1.595 39.395 1.845 40.405 ;
  LAYER M1 ;
        RECT 1.595 37.295 1.845 38.305 ;
  LAYER M1 ;
        RECT 1.165 52.415 1.415 55.945 ;
  LAYER M1 ;
        RECT 1.165 46.535 1.415 50.065 ;
  LAYER M1 ;
        RECT 1.165 40.655 1.415 44.185 ;
  LAYER M1 ;
        RECT 2.025 52.415 2.275 55.945 ;
  LAYER M1 ;
        RECT 2.025 46.535 2.275 50.065 ;
  LAYER M1 ;
        RECT 2.025 40.655 2.275 44.185 ;
  LAYER M1 ;
        RECT 2.455 52.415 2.705 55.945 ;
  LAYER M1 ;
        RECT 2.455 51.155 2.705 52.165 ;
  LAYER M1 ;
        RECT 2.455 46.535 2.705 50.065 ;
  LAYER M1 ;
        RECT 2.455 45.275 2.705 46.285 ;
  LAYER M1 ;
        RECT 2.455 40.655 2.705 44.185 ;
  LAYER M1 ;
        RECT 2.455 39.395 2.705 40.405 ;
  LAYER M1 ;
        RECT 2.455 37.295 2.705 38.305 ;
  LAYER M1 ;
        RECT 2.885 52.415 3.135 55.945 ;
  LAYER M1 ;
        RECT 2.885 46.535 3.135 50.065 ;
  LAYER M1 ;
        RECT 2.885 40.655 3.135 44.185 ;
  LAYER M1 ;
        RECT 3.315 52.415 3.565 55.945 ;
  LAYER M1 ;
        RECT 3.315 51.155 3.565 52.165 ;
  LAYER M1 ;
        RECT 3.315 46.535 3.565 50.065 ;
  LAYER M1 ;
        RECT 3.315 45.275 3.565 46.285 ;
  LAYER M1 ;
        RECT 3.315 40.655 3.565 44.185 ;
  LAYER M1 ;
        RECT 3.315 39.395 3.565 40.405 ;
  LAYER M1 ;
        RECT 3.315 37.295 3.565 38.305 ;
  LAYER M1 ;
        RECT 3.745 52.415 3.995 55.945 ;
  LAYER M1 ;
        RECT 3.745 46.535 3.995 50.065 ;
  LAYER M1 ;
        RECT 3.745 40.655 3.995 44.185 ;
  LAYER M2 ;
        RECT 1.55 55.72 3.61 56 ;
  LAYER M2 ;
        RECT 1.55 51.52 3.61 51.8 ;
  LAYER M2 ;
        RECT 1.12 55.3 4.04 55.58 ;
  LAYER M2 ;
        RECT 1.55 49.84 3.61 50.12 ;
  LAYER M2 ;
        RECT 1.55 45.64 3.61 45.92 ;
  LAYER M2 ;
        RECT 1.12 49.42 4.04 49.7 ;
  LAYER M2 ;
        RECT 1.55 43.96 3.61 44.24 ;
  LAYER M2 ;
        RECT 1.55 39.76 3.61 40.04 ;
  LAYER M2 ;
        RECT 1.12 43.54 4.04 43.82 ;
  LAYER M2 ;
        RECT 1.55 37.66 3.61 37.94 ;
  LAYER M3 ;
        RECT 2.01 43.94 2.29 56.02 ;
  LAYER M3 ;
        RECT 2.44 39.74 2.72 51.82 ;
  LAYER M3 ;
        RECT 2.87 43.52 3.15 55.6 ;
  LAYER M1 ;
        RECT 8.475 52.415 8.725 55.945 ;
  LAYER M1 ;
        RECT 8.475 51.155 8.725 52.165 ;
  LAYER M1 ;
        RECT 8.475 46.535 8.725 50.065 ;
  LAYER M1 ;
        RECT 8.475 45.275 8.725 46.285 ;
  LAYER M1 ;
        RECT 8.475 40.655 8.725 44.185 ;
  LAYER M1 ;
        RECT 8.475 39.395 8.725 40.405 ;
  LAYER M1 ;
        RECT 8.475 37.295 8.725 38.305 ;
  LAYER M1 ;
        RECT 8.905 52.415 9.155 55.945 ;
  LAYER M1 ;
        RECT 8.905 46.535 9.155 50.065 ;
  LAYER M1 ;
        RECT 8.905 40.655 9.155 44.185 ;
  LAYER M1 ;
        RECT 8.045 52.415 8.295 55.945 ;
  LAYER M1 ;
        RECT 8.045 46.535 8.295 50.065 ;
  LAYER M1 ;
        RECT 8.045 40.655 8.295 44.185 ;
  LAYER M1 ;
        RECT 7.615 52.415 7.865 55.945 ;
  LAYER M1 ;
        RECT 7.615 51.155 7.865 52.165 ;
  LAYER M1 ;
        RECT 7.615 46.535 7.865 50.065 ;
  LAYER M1 ;
        RECT 7.615 45.275 7.865 46.285 ;
  LAYER M1 ;
        RECT 7.615 40.655 7.865 44.185 ;
  LAYER M1 ;
        RECT 7.615 39.395 7.865 40.405 ;
  LAYER M1 ;
        RECT 7.615 37.295 7.865 38.305 ;
  LAYER M1 ;
        RECT 7.185 52.415 7.435 55.945 ;
  LAYER M1 ;
        RECT 7.185 46.535 7.435 50.065 ;
  LAYER M1 ;
        RECT 7.185 40.655 7.435 44.185 ;
  LAYER M1 ;
        RECT 6.755 52.415 7.005 55.945 ;
  LAYER M1 ;
        RECT 6.755 51.155 7.005 52.165 ;
  LAYER M1 ;
        RECT 6.755 46.535 7.005 50.065 ;
  LAYER M1 ;
        RECT 6.755 45.275 7.005 46.285 ;
  LAYER M1 ;
        RECT 6.755 40.655 7.005 44.185 ;
  LAYER M1 ;
        RECT 6.755 39.395 7.005 40.405 ;
  LAYER M1 ;
        RECT 6.755 37.295 7.005 38.305 ;
  LAYER M1 ;
        RECT 6.325 52.415 6.575 55.945 ;
  LAYER M1 ;
        RECT 6.325 46.535 6.575 50.065 ;
  LAYER M1 ;
        RECT 6.325 40.655 6.575 44.185 ;
  LAYER M2 ;
        RECT 6.71 55.72 8.77 56 ;
  LAYER M2 ;
        RECT 6.71 51.52 8.77 51.8 ;
  LAYER M2 ;
        RECT 6.28 55.3 9.2 55.58 ;
  LAYER M2 ;
        RECT 6.71 49.84 8.77 50.12 ;
  LAYER M2 ;
        RECT 6.71 45.64 8.77 45.92 ;
  LAYER M2 ;
        RECT 6.28 49.42 9.2 49.7 ;
  LAYER M2 ;
        RECT 6.71 43.96 8.77 44.24 ;
  LAYER M2 ;
        RECT 6.71 39.76 8.77 40.04 ;
  LAYER M2 ;
        RECT 6.28 43.54 9.2 43.82 ;
  LAYER M2 ;
        RECT 6.71 37.66 8.77 37.94 ;
  LAYER M3 ;
        RECT 8.03 43.94 8.31 56.02 ;
  LAYER M3 ;
        RECT 7.6 39.74 7.88 51.82 ;
  LAYER M3 ;
        RECT 7.17 43.52 7.45 55.6 ;
  END 
END CURRENT_MIRROR_OTA
