MACRO DCL_PMOS_S_70252776_X3_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN DCL_PMOS_S_70252776_X3_Y1 0 0 ;
  SIZE 4300 BY 7560 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 260 2290 4780 ;
    END
  END D
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2440 680 2720 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 7225 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 7225 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M2 ;
      RECT 1120 280 3180 560 ;
    LAYER M2 ;
      RECT 1120 4480 3180 4760 ;
    LAYER M2 ;
      RECT 690 700 3610 980 ;
    LAYER M2 ;
      RECT 1120 6580 3180 6860 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6635 3095 6805 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6635 2235 6805 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V2 ;
      RECT 2075 345 2225 495 ;
    LAYER V2 ;
      RECT 2075 4545 2225 4695 ;
    LAYER V2 ;
      RECT 2505 765 2655 915 ;
    LAYER V2 ;
      RECT 2505 6645 2655 6795 ;
  END
END DCL_PMOS_S_70252776_X3_Y1
