MACRO NMOS_S_89651636_X9_Y2
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_89651636_X9_Y2 0 0 ;
  SIZE 9460 BY 13440 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4160 260 4440 6460 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4590 4460 4870 10660 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5020 680 5300 12760 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 13105 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 13105 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 13105 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 13105 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 13105 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 13105 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 13105 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 13105 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 8045 335 8295 3865 ;
    LAYER M1 ;
      RECT 8045 4115 8295 5125 ;
    LAYER M1 ;
      RECT 8045 6215 8295 9745 ;
    LAYER M1 ;
      RECT 8045 9995 8295 11005 ;
    LAYER M1 ;
      RECT 8045 12095 8295 13105 ;
    LAYER M1 ;
      RECT 8475 335 8725 3865 ;
    LAYER M1 ;
      RECT 8475 6215 8725 9745 ;
    LAYER M2 ;
      RECT 1120 280 8340 560 ;
    LAYER M2 ;
      RECT 1120 4480 8340 4760 ;
    LAYER M2 ;
      RECT 690 700 8770 980 ;
    LAYER M2 ;
      RECT 1120 6160 8340 6440 ;
    LAYER M2 ;
      RECT 1120 10360 8340 10640 ;
    LAYER M2 ;
      RECT 690 6580 8770 6860 ;
    LAYER M2 ;
      RECT 1120 12460 8340 12740 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12515 1375 12685 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12515 2235 12685 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12515 3095 12685 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12515 3955 12685 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12515 4815 12685 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12515 5675 12685 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12515 6535 12685 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12515 7395 12685 ;
    LAYER V1 ;
      RECT 8085 335 8255 505 ;
    LAYER V1 ;
      RECT 8085 4535 8255 4705 ;
    LAYER V1 ;
      RECT 8085 6215 8255 6385 ;
    LAYER V1 ;
      RECT 8085 10415 8255 10585 ;
    LAYER V1 ;
      RECT 8085 12515 8255 12685 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 8515 755 8685 925 ;
    LAYER V1 ;
      RECT 8515 6635 8685 6805 ;
    LAYER V2 ;
      RECT 4225 345 4375 495 ;
    LAYER V2 ;
      RECT 4225 6225 4375 6375 ;
    LAYER V2 ;
      RECT 4655 4545 4805 4695 ;
    LAYER V2 ;
      RECT 4655 10425 4805 10575 ;
    LAYER V2 ;
      RECT 5085 765 5235 915 ;
    LAYER V2 ;
      RECT 5085 6645 5235 6795 ;
    LAYER V2 ;
      RECT 5085 12525 5235 12675 ;
  END
END NMOS_S_89651636_X9_Y2
